// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/CAPTURE_VIRTEX.v,v 1.8.22.1 2003/11/18 20:41:33 wloo Exp $
/*

FUNCTION	: Special Function Cell, CAPTURE_VIRTEX

*/

`timescale  100 ps / 10 ps


module CAPTURE_VIRTEX (CAP, CLK);

    input  CAP, CLK;

endmodule

