// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/CAPTURE_FPGACORE.v,v 1.1.20.1 2003/11/18 20:41:33 wloo Exp $
/*

FUNCTION	: Special Function Cell, CAPTURE_FPGACORE

*/

`timescale  100 ps / 10 ps


module CAPTURE_FPGACORE (CAP, CLK);

    input  CAP, CLK;

endmodule

