// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/VCC.v,v 1.8.22.1 2003/11/18 20:41:40 wloo Exp $

/*

FUNCTION	: VCC cell

*/

`timescale  100 ps / 10 ps


module VCC(P);

    output P;

	assign P = 1'b1;

endmodule

