// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/PPC405_ADV.v,v 1.1.4.7 2004/09/15 15:59:30 patrickp Exp $

`timescale 1 ps / 1 ps

module PPC405_ADV (
	APUFCMDECODED,
	APUFCMDECUDI,
	APUFCMDECUDIVALID,
	APUFCMENDIAN,
	APUFCMFLUSH,
	APUFCMINSTRUCTION,
	APUFCMINSTRVALID,
	APUFCMLOADBYTEEN,
	APUFCMLOADDATA,
	APUFCMLOADDVALID,
	APUFCMOPERANDVALID,
	APUFCMRADATA,
	APUFCMRBDATA,
	APUFCMWRITEBACKOK,
	APUFCMXERCA,
	C405CPMCORESLEEPREQ,
	C405CPMMSRCE,
	C405CPMMSREE,
	C405CPMTIMERIRQ,
	C405CPMTIMERRESETREQ,
	C405DBGLOADDATAONAPUDBUS,
	C405DBGMSRWE,
	C405DBGSTOPACK,
	C405DBGWBCOMPLETE,
	C405DBGWBFULL,
	C405DBGWBIAR,
	C405JTGCAPTUREDR,
	C405JTGEXTEST,
	C405JTGPGMOUT,
	C405JTGSHIFTDR,
	C405JTGTDO,
	C405JTGTDOEN,
	C405JTGUPDATEDR,
	C405PLBDCUABORT,
	C405PLBDCUABUS,
	C405PLBDCUBE,
	C405PLBDCUCACHEABLE,
	C405PLBDCUGUARDED,
	C405PLBDCUPRIORITY,
	C405PLBDCUREQUEST,
	C405PLBDCURNW,
	C405PLBDCUSIZE2,
	C405PLBDCUU0ATTR,
	C405PLBDCUWRDBUS,
	C405PLBDCUWRITETHRU,
	C405PLBICUABORT,
	C405PLBICUABUS,
	C405PLBICUCACHEABLE,
	C405PLBICUPRIORITY,
	C405PLBICUREQUEST,
	C405PLBICUSIZE,
	C405PLBICUU0ATTR,
	C405RSTCHIPRESETREQ,
	C405RSTCORERESETREQ,
	C405RSTSYSRESETREQ,
	C405TRCCYCLE,
	C405TRCEVENEXECUTIONSTATUS,
	C405TRCODDEXECUTIONSTATUS,
	C405TRCTRACESTATUS,
	C405TRCTRIGGEREVENTOUT,
	C405TRCTRIGGEREVENTTYPE,
	C405XXXMACHINECHECK,
	DCREMACABUS,
	DCREMACCLK,
	DCREMACDBUS,
	DCREMACENABLER,
	DCREMACREAD,
	DCREMACWRITE,
	DSOCMBRAMABUS,
	DSOCMBRAMBYTEWRITE,
	DSOCMBRAMEN,
	DSOCMBRAMWRDBUS,
	DSOCMBUSY,
	DSOCMRDADDRVALID,
	DSOCMWRADDRVALID,
	EXTDCRABUS,
	EXTDCRDBUSOUT,
	EXTDCRREAD,
	EXTDCRWRITE,
	ISOCMBRAMEN,
	ISOCMBRAMEVENWRITEEN,
	ISOCMBRAMODDWRITEEN,
	ISOCMBRAMRDABUS,
	ISOCMBRAMWRABUS,
	ISOCMBRAMWRDBUS,
	ISOCMDCRBRAMEVENEN,
	ISOCMDCRBRAMODDEN,
	ISOCMDCRBRAMRDSELECT,
	BRAMDSOCMCLK,
	BRAMDSOCMRDDBUS,
	BRAMISOCMCLK,
	BRAMISOCMDCRRDDBUS,
	BRAMISOCMRDDBUS,
	CPMC405CLOCK,
	CPMC405CORECLKINACTIVE,
	CPMC405CPUCLKEN,
	CPMC405JTAGCLKEN,
	CPMC405SYNCBYPASS,
	CPMC405TIMERCLKEN,
	CPMC405TIMERTICK,
	CPMDCRCLK,
	CPMFCMCLK,
	DBGC405DEBUGHALT,
	DBGC405EXTBUSHOLDACK,
	DBGC405UNCONDDEBUGEVENT,
	DSARCVALUE,
	DSCNTLVALUE,
	DSOCMRWCOMPLETE,
	EICC405CRITINPUTIRQ,
	EICC405EXTINPUTIRQ,
	EMACDCRACK,
	EMACDCRDBUS,
	EXTDCRACK,
	EXTDCRDBUSIN,
	FCMAPUCR,
	FCMAPUDCDCREN,
	FCMAPUDCDFORCEALIGN,
	FCMAPUDCDFORCEBESTEERING,
	FCMAPUDCDFPUOP,
	FCMAPUDCDGPRWRITE,
	FCMAPUDCDLDSTBYTE,
	FCMAPUDCDLDSTDW,
	FCMAPUDCDLDSTHW,
	FCMAPUDCDLDSTQW,
	FCMAPUDCDLDSTWD,
	FCMAPUDCDLOAD,
	FCMAPUDCDPRIVOP,
	FCMAPUDCDRAEN,
	FCMAPUDCDRBEN,
	FCMAPUDCDSTORE,
	FCMAPUDCDTRAPBE,
	FCMAPUDCDTRAPLE,
	FCMAPUDCDUPDATE,
	FCMAPUDCDXERCAEN,
	FCMAPUDCDXEROVEN,
	FCMAPUDECODEBUSY,
	FCMAPUDONE,
	FCMAPUEXCEPTION,
	FCMAPUEXEBLOCKINGMCO,
	FCMAPUEXECRFIELD,
	FCMAPUEXENONBLOCKINGMCO,
	FCMAPUINSTRACK,
	FCMAPULOADWAIT,
	FCMAPURESULT,
	FCMAPURESULTVALID,
	FCMAPUSLEEPNOTREADY,
	FCMAPUXERCA,
	FCMAPUXEROV,
	ISARCVALUE,
	ISCNTLVALUE,
	JTGC405BNDSCANTDO,
	JTGC405TCK,
	JTGC405TDI,
	JTGC405TMS,
	JTGC405TRSTNEG,
	MCBCPUCLKEN,
	MCBJTAGEN,
	MCBTIMEREN,
	MCPPCRST,
	PLBC405DCUADDRACK,
	PLBC405DCUBUSY,
	PLBC405DCUERR,
	PLBC405DCURDDACK,
	PLBC405DCURDDBUS,
	PLBC405DCURDWDADDR,
	PLBC405DCUSSIZE1,
	PLBC405DCUWRDACK,
	PLBC405ICUADDRACK,
	PLBC405ICUBUSY,
	PLBC405ICUERR,
	PLBC405ICURDDACK,
	PLBC405ICURDDBUS,
	PLBC405ICURDWDADDR,
	PLBC405ICUSSIZE1,
	PLBCLK,
	RSTC405RESETCHIP,
	RSTC405RESETCORE,
	RSTC405RESETSYS,
	TIEAPUCONTROL,
	TIEAPUUDI1,
	TIEAPUUDI2,
	TIEAPUUDI3,
	TIEAPUUDI4,
	TIEAPUUDI5,
	TIEAPUUDI6,
	TIEAPUUDI7,
	TIEAPUUDI8,
	TIEC405DETERMINISTICMULT,
	TIEC405DISOPERANDFWD,
	TIEC405MMUEN,
	TIEDCRADDR,
	TIEPVRBIT10,
	TIEPVRBIT11,
	TIEPVRBIT28,
	TIEPVRBIT29,
	TIEPVRBIT30,
	TIEPVRBIT31,
	TIEPVRBIT8,
	TIEPVRBIT9,
	TRCC405TRACEDISABLE,
	TRCC405TRIGGEREVENTIN
);

parameter in_delay=100;
parameter out_delay=100;

output APUFCMDECODED;
output APUFCMDECUDIVALID;
output APUFCMENDIAN;
output APUFCMFLUSH;
output APUFCMINSTRVALID;
output APUFCMLOADDVALID;
output APUFCMOPERANDVALID;
output APUFCMWRITEBACKOK;
output APUFCMXERCA;
output C405CPMCORESLEEPREQ;
output C405CPMMSRCE;
output C405CPMMSREE;
output C405CPMTIMERIRQ;
output C405CPMTIMERRESETREQ;
output C405DBGLOADDATAONAPUDBUS;
output C405DBGMSRWE;
output C405DBGSTOPACK;
output C405DBGWBCOMPLETE;
output C405DBGWBFULL;
output C405JTGCAPTUREDR;
output C405JTGEXTEST;
output C405JTGPGMOUT;
output C405JTGSHIFTDR;
output C405JTGTDO;
output C405JTGTDOEN;
output C405JTGUPDATEDR;
output C405PLBDCUABORT;
output C405PLBDCUCACHEABLE;
output C405PLBDCUGUARDED;
output C405PLBDCUREQUEST;
output C405PLBDCURNW;
output C405PLBDCUSIZE2;
output C405PLBDCUU0ATTR;
output C405PLBDCUWRITETHRU;
output C405PLBICUABORT;
output C405PLBICUCACHEABLE;
output C405PLBICUREQUEST;
output C405PLBICUU0ATTR;
output C405RSTCHIPRESETREQ;
output C405RSTCORERESETREQ;
output C405RSTSYSRESETREQ;
output C405TRCCYCLE;
output C405TRCTRIGGEREVENTOUT;
output C405XXXMACHINECHECK;
output DCREMACCLK;
output DCREMACENABLER;
output DCREMACREAD;
output DCREMACWRITE;
output DSOCMBRAMEN;
output DSOCMBUSY;
output DSOCMRDADDRVALID;
output DSOCMWRADDRVALID;
output EXTDCRREAD;
output EXTDCRWRITE;
output ISOCMBRAMEN;
output ISOCMBRAMEVENWRITEEN;
output ISOCMBRAMODDWRITEEN;
output ISOCMDCRBRAMEVENEN;
output ISOCMDCRBRAMODDEN;
output ISOCMDCRBRAMRDSELECT;
output [0:10] C405TRCTRIGGEREVENTTYPE;
output [0:1] C405PLBDCUPRIORITY;
output [0:1] C405PLBICUPRIORITY;
output [0:1] C405TRCEVENEXECUTIONSTATUS;
output [0:1] C405TRCODDEXECUTIONSTATUS;
output [0:29] C405DBGWBIAR;
output [0:29] C405PLBICUABUS;
output [0:2] APUFCMDECUDI;
output [0:31] APUFCMINSTRUCTION;
output [0:31] APUFCMLOADDATA;
output [0:31] APUFCMRADATA;
output [0:31] APUFCMRBDATA;
output [0:31] C405PLBDCUABUS;
output [0:31] DCREMACDBUS;
output [0:31] DSOCMBRAMWRDBUS;
output [0:31] EXTDCRDBUSOUT;
output [0:31] ISOCMBRAMWRDBUS;
output [0:3] APUFCMLOADBYTEEN;
output [0:3] C405TRCTRACESTATUS;
output [0:3] DSOCMBRAMBYTEWRITE;
output [0:63] C405PLBDCUWRDBUS;
output [0:7] C405PLBDCUBE;
output [0:9] EXTDCRABUS;
output [2:3] C405PLBICUSIZE;
output [8:28] ISOCMBRAMRDABUS;
output [8:28] ISOCMBRAMWRABUS;
output [8:29] DSOCMBRAMABUS;
output [8:9] DCREMACABUS;

input BRAMDSOCMCLK;
input BRAMISOCMCLK;
input CPMC405CLOCK;
input CPMC405CORECLKINACTIVE;
input CPMC405CPUCLKEN;
input CPMC405JTAGCLKEN;
input CPMC405SYNCBYPASS;
input CPMC405TIMERCLKEN;
input CPMC405TIMERTICK;
input CPMDCRCLK;
input CPMFCMCLK;
input DBGC405DEBUGHALT;
input DBGC405EXTBUSHOLDACK;
input DBGC405UNCONDDEBUGEVENT;
input DSOCMRWCOMPLETE;
input EICC405CRITINPUTIRQ;
input EICC405EXTINPUTIRQ;
input EMACDCRACK;
input EXTDCRACK;
input FCMAPUDCDCREN;
input FCMAPUDCDFORCEALIGN;
input FCMAPUDCDFORCEBESTEERING;
input FCMAPUDCDFPUOP;
input FCMAPUDCDGPRWRITE;
input FCMAPUDCDLDSTBYTE;
input FCMAPUDCDLDSTDW;
input FCMAPUDCDLDSTHW;
input FCMAPUDCDLDSTQW;
input FCMAPUDCDLDSTWD;
input FCMAPUDCDLOAD;
input FCMAPUDCDPRIVOP;
input FCMAPUDCDRAEN;
input FCMAPUDCDRBEN;
input FCMAPUDCDSTORE;
input FCMAPUDCDTRAPBE;
input FCMAPUDCDTRAPLE;
input FCMAPUDCDUPDATE;
input FCMAPUDCDXERCAEN;
input FCMAPUDCDXEROVEN;
input FCMAPUDECODEBUSY;
input FCMAPUDONE;
input FCMAPUEXCEPTION;
input FCMAPUEXEBLOCKINGMCO;
input FCMAPUEXENONBLOCKINGMCO;
input FCMAPUINSTRACK;
input FCMAPULOADWAIT;
input FCMAPURESULTVALID;
input FCMAPUSLEEPNOTREADY;
input FCMAPUXERCA;
input FCMAPUXEROV;
input JTGC405BNDSCANTDO;
input JTGC405TCK;
input JTGC405TDI;
input JTGC405TMS;
input JTGC405TRSTNEG;
input MCBCPUCLKEN;
input MCBJTAGEN;
input MCBTIMEREN;
input MCPPCRST;
input PLBC405DCUADDRACK;
input PLBC405DCUBUSY;
input PLBC405DCUERR;
input PLBC405DCURDDACK;
input PLBC405DCUSSIZE1;
input PLBC405DCUWRDACK;
input PLBC405ICUADDRACK;
input PLBC405ICUBUSY;
input PLBC405ICUERR;
input PLBC405ICURDDACK;
input PLBC405ICUSSIZE1;
input PLBCLK;
input RSTC405RESETCHIP;
input RSTC405RESETCORE;
input RSTC405RESETSYS;
input TIEC405DETERMINISTICMULT;
input TIEC405DISOPERANDFWD;
input TIEC405MMUEN;
input TIEPVRBIT10;
input TIEPVRBIT11;
input TIEPVRBIT28;
input TIEPVRBIT29;
input TIEPVRBIT30;
input TIEPVRBIT31;
input TIEPVRBIT8;
input TIEPVRBIT9;
input TRCC405TRACEDISABLE;
input TRCC405TRIGGEREVENTIN;
input [0:15] TIEAPUCONTROL;
input [0:23] TIEAPUUDI1;
input [0:23] TIEAPUUDI2;
input [0:23] TIEAPUUDI3;
input [0:23] TIEAPUUDI4;
input [0:23] TIEAPUUDI5;
input [0:23] TIEAPUUDI6;
input [0:23] TIEAPUUDI7;
input [0:23] TIEAPUUDI8;
input [0:2] FCMAPUEXECRFIELD;
input [0:31] BRAMDSOCMRDDBUS;
input [0:31] BRAMISOCMDCRRDDBUS;
input [0:31] EMACDCRDBUS;
input [0:31] EXTDCRDBUSIN;
input [0:31] FCMAPURESULT;
input [0:3] FCMAPUCR;
input [0:5] TIEDCRADDR;
input [0:63] BRAMISOCMRDDBUS;
input [0:63] PLBC405DCURDDBUS;
input [0:63] PLBC405ICURDDBUS;
input [0:7] DSARCVALUE;
input [0:7] DSCNTLVALUE;
input [0:7] ISARCVALUE;
input [0:7] ISCNTLVALUE;
input [1:3] PLBC405DCURDWDADDR;
input [1:3] PLBC405ICURDWDADDR;

wire APUFCMDECODED_delay;
wire APUFCMDECUDIVALID_delay;
wire APUFCMENDIAN_delay;
wire APUFCMFLUSH_delay;
wire APUFCMINSTRVALID_delay;
wire APUFCMLOADDVALID_delay;
wire APUFCMOPERANDVALID_delay;
wire APUFCMWRITEBACKOK_delay;
wire APUFCMXERCA_delay;
wire BRAMDSOCMCLK_delay;
wire BRAMISOCMCLK_delay;
wire C405CPMCORESLEEPREQ_delay;
wire C405CPMMSRCE_delay;
wire C405CPMMSREE_delay;
wire C405CPMTIMERIRQ_delay;
wire C405CPMTIMERRESETREQ_delay;
wire C405DBGLOADDATAONAPUDBUS_delay;
wire C405DBGMSRWE_delay;
wire C405DBGSTOPACK_delay;
wire C405DBGWBCOMPLETE_delay;
wire C405DBGWBFULL_delay;
wire C405JTGCAPTUREDR_delay;
wire C405JTGEXTEST_delay;
wire C405JTGPGMOUT_delay;
wire C405JTGSHIFTDR_delay;
wire C405JTGTDOEN_delay;
wire C405JTGTDO_delay;
wire C405JTGUPDATEDR_delay;
wire C405PLBDCUABORT_delay;
wire C405PLBDCUCACHEABLE_delay;
wire C405PLBDCUGUARDED_delay;
wire C405PLBDCUREQUEST_delay;
wire C405PLBDCURNW_delay;
wire C405PLBDCUSIZE2_delay;
wire C405PLBDCUU0ATTR_delay;
wire C405PLBDCUWRITETHRU_delay;
wire C405PLBICUABORT_delay;
wire C405PLBICUCACHEABLE_delay;
wire C405PLBICUREQUEST_delay;
wire C405PLBICUU0ATTR_delay;
wire C405RSTCHIPRESETREQ_delay;
wire C405RSTCORERESETREQ_delay;
wire C405RSTSYSRESETREQ_delay;
wire C405TRCCYCLE_delay;
wire C405TRCTRIGGEREVENTOUT_delay;
wire C405XXXMACHINECHECK_delay;
wire CPMC405CLOCK_delay;
wire CPMC405CORECLKINACTIVE_delay;
wire CPMC405CPUCLKEN_delay;
wire CPMC405JTAGCLKEN_delay;
wire CPMC405SYNCBYPASS_delay;
wire CPMC405TIMERCLKEN_delay;
wire CPMC405TIMERTICK_delay;
wire CPMDCRCLK_delay;
wire CPMFCMCLK_delay;
wire DBGC405DEBUGHALT_delay;
wire DBGC405EXTBUSHOLDACK_delay;
wire DBGC405UNCONDDEBUGEVENT_delay;
wire DCREMACCLK_delay;
wire DCREMACENABLER_delay;
wire DCREMACREAD_delay;
wire DCREMACWRITE_delay;
wire DSOCMBRAMEN_delay;
wire DSOCMBUSY_delay;
wire DSOCMRDADDRVALID_delay;
wire DSOCMRWCOMPLETE_delay;
wire DSOCMWRADDRVALID_delay;
wire EICC405CRITINPUTIRQ_delay;
wire EICC405EXTINPUTIRQ_delay;
wire EMACDCRACK_delay;
wire EXTDCRACK_delay;
wire EXTDCRREAD_delay;
wire EXTDCRWRITE_delay;
wire FCMAPUDCDCREN_delay;
wire FCMAPUDCDFORCEALIGN_delay;
wire FCMAPUDCDFORCEBESTEERING_delay;
wire FCMAPUDCDFPUOP_delay;
wire FCMAPUDCDGPRWRITE_delay;
wire FCMAPUDCDLDSTBYTE_delay;
wire FCMAPUDCDLDSTDW_delay;
wire FCMAPUDCDLDSTHW_delay;
wire FCMAPUDCDLDSTQW_delay;
wire FCMAPUDCDLDSTWD_delay;
wire FCMAPUDCDLOAD_delay;
wire FCMAPUDCDPRIVOP_delay;
wire FCMAPUDCDRAEN_delay;
wire FCMAPUDCDRBEN_delay;
wire FCMAPUDCDSTORE_delay;
wire FCMAPUDCDTRAPBE_delay;
wire FCMAPUDCDTRAPLE_delay;
wire FCMAPUDCDUPDATE_delay;
wire FCMAPUDCDXERCAEN_delay;
wire FCMAPUDCDXEROVEN_delay;
wire FCMAPUDECODEBUSY_delay;
wire FCMAPUDONE_delay;
wire FCMAPUEXCEPTION_delay;
wire FCMAPUEXEBLOCKINGMCO_delay;
wire FCMAPUEXENONBLOCKINGMCO_delay;
wire FCMAPUINSTRACK_delay;
wire FCMAPULOADWAIT_delay;
wire FCMAPURESULTVALID_delay;
wire FCMAPUSLEEPNOTREADY_delay;
wire FCMAPUXERCA_delay;
wire FCMAPUXEROV_delay;
wire ISOCMBRAMEN_delay;
wire ISOCMBRAMEVENWRITEEN_delay;
wire ISOCMBRAMODDWRITEEN_delay;
wire ISOCMDCRBRAMEVENEN_delay;
wire ISOCMDCRBRAMODDEN_delay;
wire ISOCMDCRBRAMRDSELECT_delay;
wire JTGC405BNDSCANTDO_delay;
wire JTGC405TCK_delay;
wire JTGC405TDI_delay;
wire JTGC405TMS_delay;
wire JTGC405TRSTNEG_delay;
wire MCBCPUCLKEN_delay;
wire MCBJTAGEN_delay;
wire MCBTIMEREN_delay;
wire MCPPCRST_delay;
wire PLBC405DCUADDRACK_delay;
wire PLBC405DCUBUSY_delay;
wire PLBC405DCUERR_delay;
wire PLBC405DCURDDACK_delay;
wire PLBC405DCUSSIZE1_delay;
wire PLBC405DCUWRDACK_delay;
wire PLBC405ICUADDRACK_delay;
wire PLBC405ICUBUSY_delay;
wire PLBC405ICUERR_delay;
wire PLBC405ICURDDACK_delay;
wire PLBC405ICUSSIZE1_delay;
wire PLBCLK_delay;
wire RSTC405RESETCHIP_delay;
wire RSTC405RESETCORE_delay;
wire RSTC405RESETSYS_delay;
wire TIEC405DETERMINISTICMULT_delay;
wire TIEC405DISOPERANDFWD_delay;
wire TIEC405MMUEN_delay;
wire TIEPVRBIT10_delay;
wire TIEPVRBIT11_delay;
wire TIEPVRBIT28_delay;
wire TIEPVRBIT29_delay;
wire TIEPVRBIT30_delay;
wire TIEPVRBIT31_delay;
wire TIEPVRBIT8_delay;
wire TIEPVRBIT9_delay;
wire TRCC405TRACEDISABLE_delay;
wire TRCC405TRIGGEREVENTIN_delay;
wire [0:10] C405TRCTRIGGEREVENTTYPE_delay;
wire [0:15] TIEAPUCONTROL_delay;
wire [0:1] C405PLBDCUPRIORITY_delay;
wire [0:1] C405PLBICUPRIORITY_delay;
wire [0:1] C405TRCEVENEXECUTIONSTATUS_delay;
wire [0:1] C405TRCODDEXECUTIONSTATUS_delay;
wire [0:23] TIEAPUUDI1_delay;
wire [0:23] TIEAPUUDI2_delay;
wire [0:23] TIEAPUUDI3_delay;
wire [0:23] TIEAPUUDI4_delay;
wire [0:23] TIEAPUUDI5_delay;
wire [0:23] TIEAPUUDI6_delay;
wire [0:23] TIEAPUUDI7_delay;
wire [0:23] TIEAPUUDI8_delay;
wire [0:29] C405DBGWBIAR_delay;
wire [0:29] C405PLBICUABUS_delay;
wire [0:2] APUFCMDECUDI_delay;
wire [0:2] FCMAPUEXECRFIELD_delay;
wire [0:31] APUFCMINSTRUCTION_delay;
wire [0:31] APUFCMLOADDATA_delay;
wire [0:31] APUFCMRADATA_delay;
wire [0:31] APUFCMRBDATA_delay;
wire [0:31] BRAMDSOCMRDDBUS_delay;
wire [0:31] BRAMISOCMDCRRDDBUS_delay;
wire [0:31] C405PLBDCUABUS_delay;
wire [0:31] DCREMACDBUS_delay;
wire [0:31] DSOCMBRAMWRDBUS_delay;
wire [0:31] EMACDCRDBUS_delay;
wire [0:31] EXTDCRDBUSIN_delay;
wire [0:31] EXTDCRDBUSOUT_delay;
wire [0:31] FCMAPURESULT_delay;
wire [0:31] ISOCMBRAMWRDBUS_delay;
wire [0:3] APUFCMLOADBYTEEN_delay;
wire [0:3] C405TRCTRACESTATUS_delay;
wire [0:3] DSOCMBRAMBYTEWRITE_delay;
wire [0:3] FCMAPUCR_delay;
wire [0:5] TIEDCRADDR_delay;
wire [0:63] BRAMISOCMRDDBUS_delay;
wire [0:63] C405PLBDCUWRDBUS_delay;
wire [0:63] PLBC405DCURDDBUS_delay;
wire [0:63] PLBC405ICURDDBUS_delay;
wire [0:7] C405PLBDCUBE_delay;
wire [0:7] DSARCVALUE_delay;
wire [0:7] DSCNTLVALUE_delay;
wire [0:7] ISARCVALUE_delay;
wire [0:7] ISCNTLVALUE_delay;
wire [0:9] EXTDCRABUS_delay;
wire [1:3] PLBC405DCURDWDADDR_delay;
wire [1:3] PLBC405ICURDWDADDR_delay;
wire [2:3] C405PLBICUSIZE_delay;
wire [8:28] ISOCMBRAMRDABUS_delay;
wire [8:28] ISOCMBRAMWRABUS_delay;
wire [8:29] DSOCMBRAMABUS_delay;
wire [8:9] DCREMACABUS_delay;

assign #(in_delay) EMACDCRACK_delay = EMACDCRACK;

assign #(in_delay) EMACDCRDBUS_delay[0:31] = EMACDCRDBUS[0:31];
assign #(in_delay) BRAMDSOCMRDDBUS_delay[0:31] = BRAMDSOCMRDDBUS[0:31];
assign #(in_delay) DSOCMRWCOMPLETE_delay = DSOCMRWCOMPLETE;
assign #(in_delay) BRAMISOCMRDDBUS_delay[0:63] = BRAMISOCMRDDBUS[0:63];
assign #(in_delay) BRAMISOCMDCRRDDBUS_delay[0:31] = BRAMISOCMDCRRDDBUS[0:31];
assign #(in_delay) CPMC405CORECLKINACTIVE_delay = CPMC405CORECLKINACTIVE;
assign #(in_delay) CPMC405CPUCLKEN_delay = CPMC405CPUCLKEN;
assign #(in_delay) CPMC405JTAGCLKEN_delay = CPMC405JTAGCLKEN;
assign #(in_delay) CPMC405TIMERCLKEN_delay = CPMC405TIMERCLKEN;
assign #(in_delay) CPMC405SYNCBYPASS_delay = CPMC405SYNCBYPASS;
assign #(in_delay) CPMC405TIMERTICK_delay = CPMC405TIMERTICK;
assign #(in_delay) DBGC405DEBUGHALT_delay = DBGC405DEBUGHALT;
assign #(in_delay) DBGC405EXTBUSHOLDACK_delay = DBGC405EXTBUSHOLDACK;
assign #(in_delay) DBGC405UNCONDDEBUGEVENT_delay = DBGC405UNCONDDEBUGEVENT;
assign #(in_delay) EXTDCRACK_delay = EXTDCRACK;
assign #(in_delay) EXTDCRDBUSIN_delay[0:31] = EXTDCRDBUSIN[0:31];
assign #(in_delay) DSARCVALUE_delay[0:7] = DSARCVALUE[0:7];
assign #(in_delay) DSCNTLVALUE_delay[0:7] = DSCNTLVALUE[0:7];
assign #(in_delay) EICC405CRITINPUTIRQ_delay = EICC405CRITINPUTIRQ;
assign #(in_delay) EICC405EXTINPUTIRQ_delay = EICC405EXTINPUTIRQ;
assign #(in_delay) ISARCVALUE_delay[0:7] = ISARCVALUE[0:7];
assign #(in_delay) ISCNTLVALUE_delay[0:7] = ISCNTLVALUE[0:7];
assign #(in_delay) JTGC405BNDSCANTDO_delay = JTGC405BNDSCANTDO;
assign #(in_delay) JTGC405TCK_delay = JTGC405TCK;
assign #(in_delay) JTGC405TDI_delay = JTGC405TDI;
assign #(in_delay) JTGC405TMS_delay = JTGC405TMS;
assign #(in_delay) JTGC405TRSTNEG_delay = JTGC405TRSTNEG;
assign #(in_delay) MCBCPUCLKEN_delay = MCBCPUCLKEN;
assign #(in_delay) MCBJTAGEN_delay = MCBJTAGEN;
assign #(in_delay) MCBTIMEREN_delay = MCBTIMEREN;
assign #(in_delay) MCPPCRST_delay = MCPPCRST;
assign #(in_delay) PLBC405DCUADDRACK_delay = PLBC405DCUADDRACK;
assign #(in_delay) PLBC405DCUBUSY_delay = PLBC405DCUBUSY;
assign #(in_delay) PLBC405DCUERR_delay = PLBC405DCUERR;
assign #(in_delay) PLBC405DCURDDACK_delay = PLBC405DCURDDACK;
assign #(in_delay) PLBC405DCURDDBUS_delay[0:63] = PLBC405DCURDDBUS[0:63];
assign #(in_delay) PLBC405DCURDWDADDR_delay[1:3] = PLBC405DCURDWDADDR[1:3];
assign #(in_delay) PLBC405DCUSSIZE1_delay = PLBC405DCUSSIZE1;
assign #(in_delay) PLBC405DCUWRDACK_delay = PLBC405DCUWRDACK;
assign #(in_delay) PLBC405ICUADDRACK_delay = PLBC405ICUADDRACK;
assign #(in_delay) PLBC405ICUBUSY_delay = PLBC405ICUBUSY;
assign #(in_delay) PLBC405ICUERR_delay = PLBC405ICUERR;
assign #(in_delay) PLBC405ICURDDACK_delay = PLBC405ICURDDACK;
assign #(in_delay) PLBC405ICURDDBUS_delay[0:63] = PLBC405ICURDDBUS[0:63];
assign #(in_delay) PLBC405ICURDWDADDR_delay[1:3] = PLBC405ICURDWDADDR[1:3];
assign #(in_delay) PLBC405ICUSSIZE1_delay = PLBC405ICUSSIZE1;
assign #(in_delay) RSTC405RESETCHIP_delay = RSTC405RESETCHIP;
assign #(in_delay) RSTC405RESETCORE_delay = RSTC405RESETCORE;
assign #(in_delay) RSTC405RESETSYS_delay = RSTC405RESETSYS;
assign #(in_delay) TIEC405DETERMINISTICMULT_delay = TIEC405DETERMINISTICMULT;
assign #(in_delay) TIEC405DISOPERANDFWD_delay = TIEC405DISOPERANDFWD;
assign #(in_delay) TIEC405MMUEN_delay = TIEC405MMUEN;
assign #(in_delay) TIEDCRADDR_delay[0:5] = TIEDCRADDR[0:5];
assign #(in_delay) TRCC405TRACEDISABLE_delay = TRCC405TRACEDISABLE;
assign #(in_delay) TRCC405TRIGGEREVENTIN_delay = TRCC405TRIGGEREVENTIN;
assign #(in_delay) FCMAPURESULT_delay[0:31] = FCMAPURESULT[0:31];
assign #(in_delay) FCMAPUCR_delay[0:3] = FCMAPUCR[0:3];
assign #(in_delay) FCMAPUEXECRFIELD_delay[0:2] = FCMAPUEXECRFIELD[0:2];
assign #(in_delay) FCMAPUDONE_delay = FCMAPUDONE;
assign #(in_delay) FCMAPURESULTVALID_delay = FCMAPURESULTVALID;
assign #(in_delay) FCMAPUINSTRACK_delay = FCMAPUINSTRACK;
assign #(in_delay) FCMAPUEXCEPTION_delay = FCMAPUEXCEPTION;
assign #(in_delay) FCMAPUXERCA_delay = FCMAPUXERCA;
assign #(in_delay) FCMAPUXEROV_delay = FCMAPUXEROV;
assign #(in_delay) FCMAPUDCDFPUOP_delay = FCMAPUDCDFPUOP;
assign #(in_delay) FCMAPUDCDGPRWRITE_delay = FCMAPUDCDGPRWRITE;
assign #(in_delay) FCMAPUDCDRAEN_delay = FCMAPUDCDRAEN;
assign #(in_delay) FCMAPUDCDRBEN_delay = FCMAPUDCDRBEN;
assign #(in_delay) FCMAPUDCDLOAD_delay = FCMAPUDCDLOAD;
assign #(in_delay) FCMAPUDCDSTORE_delay = FCMAPUDCDSTORE;
assign #(in_delay) FCMAPUDCDXERCAEN_delay = FCMAPUDCDXERCAEN;
assign #(in_delay) FCMAPUDCDXEROVEN_delay = FCMAPUDCDXEROVEN;
assign #(in_delay) FCMAPUDCDPRIVOP_delay = FCMAPUDCDPRIVOP;
assign #(in_delay) FCMAPUDCDCREN_delay = FCMAPUDCDCREN;
assign #(in_delay) FCMAPUDCDUPDATE_delay = FCMAPUDCDUPDATE;
assign #(in_delay) FCMAPUDCDFORCEALIGN_delay = FCMAPUDCDFORCEALIGN;
assign #(in_delay) FCMAPUDCDFORCEBESTEERING_delay = FCMAPUDCDFORCEBESTEERING;
assign #(in_delay) FCMAPUDCDLDSTBYTE_delay = FCMAPUDCDLDSTBYTE;
assign #(in_delay) FCMAPUDCDLDSTHW_delay = FCMAPUDCDLDSTHW;
assign #(in_delay) FCMAPUDCDLDSTWD_delay = FCMAPUDCDLDSTWD;
assign #(in_delay) FCMAPUDCDLDSTDW_delay = FCMAPUDCDLDSTDW;
assign #(in_delay) FCMAPUDCDLDSTQW_delay = FCMAPUDCDLDSTQW;
assign #(in_delay) FCMAPUDCDTRAPBE_delay = FCMAPUDCDTRAPBE;
assign #(in_delay) FCMAPUDCDTRAPLE_delay = FCMAPUDCDTRAPLE;
assign #(in_delay) FCMAPUEXEBLOCKINGMCO_delay = FCMAPUEXEBLOCKINGMCO;
assign #(in_delay) FCMAPUEXENONBLOCKINGMCO_delay = FCMAPUEXENONBLOCKINGMCO;
assign #(in_delay) FCMAPUSLEEPNOTREADY_delay = FCMAPUSLEEPNOTREADY;
assign #(in_delay) FCMAPULOADWAIT_delay = FCMAPULOADWAIT;
assign #(in_delay) FCMAPUDECODEBUSY_delay = FCMAPUDECODEBUSY;
assign #(in_delay) TIEAPUCONTROL_delay[0:15] = TIEAPUCONTROL[0:15];
assign #(in_delay) TIEAPUUDI1_delay[0:23] = TIEAPUUDI1[0:23];
assign #(in_delay) TIEAPUUDI2_delay[0:23] = TIEAPUUDI2[0:23];
assign #(in_delay) TIEAPUUDI3_delay[0:23] = TIEAPUUDI3[0:23];
assign #(in_delay) TIEAPUUDI4_delay[0:23] = TIEAPUUDI4[0:23];
assign #(in_delay) TIEAPUUDI5_delay[0:23] = TIEAPUUDI5[0:23];
assign #(in_delay) TIEAPUUDI6_delay[0:23] = TIEAPUUDI6[0:23];
assign #(in_delay) TIEAPUUDI7_delay[0:23] = TIEAPUUDI7[0:23];
assign #(in_delay) TIEAPUUDI8_delay[0:23] = TIEAPUUDI8[0:23];

assign #(out_delay) C405CPMCORESLEEPREQ = C405CPMCORESLEEPREQ_delay;
assign #(out_delay) C405CPMMSRCE = C405CPMMSRCE_delay;
assign #(out_delay) C405CPMMSREE = C405CPMMSREE_delay;
assign #(out_delay) C405CPMTIMERIRQ = C405CPMTIMERIRQ_delay;
assign #(out_delay) C405CPMTIMERRESETREQ = C405CPMTIMERRESETREQ_delay;
assign #(out_delay) C405DBGMSRWE = C405DBGMSRWE_delay;
assign #(out_delay) C405DBGSTOPACK = C405DBGSTOPACK_delay;
assign #(out_delay) C405DBGWBCOMPLETE = C405DBGWBCOMPLETE_delay;
assign #(out_delay) C405DBGWBFULL = C405DBGWBFULL_delay;
assign #(out_delay) C405DBGWBIAR[0:29] = C405DBGWBIAR_delay[0:29];
assign #(out_delay) EXTDCRABUS[0:9] = EXTDCRABUS_delay[0:9];
assign #(out_delay) EXTDCRDBUSOUT[0:31] = EXTDCRDBUSOUT_delay[0:31];
assign #(out_delay) DCREMACDBUS[0:31] = DCREMACDBUS_delay[0:31];
assign #(out_delay) DCREMACABUS[8:9] = DCREMACABUS_delay[8:9];
assign #(out_delay) DCREMACWRITE = DCREMACWRITE_delay;
assign #(out_delay) DCREMACREAD = DCREMACREAD_delay;
assign #(out_delay) EXTDCRREAD = EXTDCRREAD_delay;
assign #(out_delay) EXTDCRWRITE = EXTDCRWRITE_delay;
assign #(out_delay) C405JTGCAPTUREDR = C405JTGCAPTUREDR_delay;
assign #(out_delay) C405JTGEXTEST = C405JTGEXTEST_delay;
assign #(out_delay) C405JTGPGMOUT = C405JTGPGMOUT_delay;
assign #(out_delay) C405JTGSHIFTDR = C405JTGSHIFTDR_delay;
assign #(out_delay) C405JTGTDO = C405JTGTDO_delay;
assign #(out_delay) C405JTGTDOEN = C405JTGTDOEN_delay;
assign #(out_delay) C405JTGUPDATEDR = C405JTGUPDATEDR_delay;
assign #(out_delay) C405PLBDCUABORT = C405PLBDCUABORT_delay;
assign #(out_delay) C405PLBDCUABUS[0:31] = C405PLBDCUABUS_delay[0:31];
assign #(out_delay) C405PLBDCUBE[0:7] = C405PLBDCUBE_delay[0:7];
assign #(out_delay) C405PLBDCUCACHEABLE = C405PLBDCUCACHEABLE_delay;
assign #(out_delay) C405PLBDCUGUARDED = C405PLBDCUGUARDED_delay;
assign #(out_delay) C405PLBDCUPRIORITY[0:1] = C405PLBDCUPRIORITY_delay[0:1];
assign #(out_delay) C405PLBDCUREQUEST = C405PLBDCUREQUEST_delay;
assign #(out_delay) C405PLBDCURNW = C405PLBDCURNW_delay;
assign #(out_delay) C405PLBDCUSIZE2 = C405PLBDCUSIZE2_delay;
assign #(out_delay) C405PLBDCUU0ATTR = C405PLBDCUU0ATTR_delay;
assign #(out_delay) C405PLBDCUWRDBUS[0:63] = C405PLBDCUWRDBUS_delay[0:63];
assign #(out_delay) C405PLBDCUWRITETHRU = C405PLBDCUWRITETHRU_delay;
assign #(out_delay) C405PLBICUABORT = C405PLBICUABORT_delay;
assign #(out_delay) C405PLBICUABUS[0:29] = C405PLBICUABUS_delay[0:29];
assign #(out_delay) C405PLBICUCACHEABLE = C405PLBICUCACHEABLE_delay;
assign #(out_delay) C405PLBICUPRIORITY[0:1] = C405PLBICUPRIORITY_delay[0:1];
assign #(out_delay) C405PLBICUREQUEST = C405PLBICUREQUEST_delay;
assign #(out_delay) C405PLBICUSIZE[2:3] = C405PLBICUSIZE_delay[2:3];
assign #(out_delay) C405PLBICUU0ATTR = C405PLBICUU0ATTR_delay;
assign #(out_delay) C405RSTCHIPRESETREQ = C405RSTCHIPRESETREQ_delay;
assign #(out_delay) C405RSTCORERESETREQ = C405RSTCORERESETREQ_delay;
assign #(out_delay) C405RSTSYSRESETREQ = C405RSTSYSRESETREQ_delay;
assign #(out_delay) C405TRCCYCLE = C405TRCCYCLE_delay;
assign #(out_delay) C405TRCEVENEXECUTIONSTATUS[0:1] = C405TRCEVENEXECUTIONSTATUS_delay[0:1];
assign #(out_delay) C405TRCODDEXECUTIONSTATUS[0:1] = C405TRCODDEXECUTIONSTATUS_delay[0:1];
assign #(out_delay) C405TRCTRACESTATUS[0:3] = C405TRCTRACESTATUS_delay[0:3];
assign #(out_delay) C405TRCTRIGGEREVENTOUT = C405TRCTRIGGEREVENTOUT_delay;
assign #(out_delay) C405TRCTRIGGEREVENTTYPE[0:10] = C405TRCTRIGGEREVENTTYPE_delay[0:10];
assign #(out_delay) C405XXXMACHINECHECK = C405XXXMACHINECHECK_delay;
assign #(out_delay) DCREMACENABLER = DCREMACENABLER_delay;
assign #(out_delay) DSOCMBRAMABUS[8:29] = DSOCMBRAMABUS_delay[8:29];
assign #(out_delay) DSOCMBRAMBYTEWRITE[0:3] = DSOCMBRAMBYTEWRITE_delay[0:3];
assign #(out_delay) DSOCMBRAMEN = DSOCMBRAMEN_delay;
assign #(out_delay) DSOCMBRAMWRDBUS[0:31] = DSOCMBRAMWRDBUS_delay[0:31];
assign #(out_delay) DSOCMBUSY = DSOCMBUSY_delay;
assign #(out_delay) DSOCMWRADDRVALID = DSOCMWRADDRVALID_delay;
assign #(out_delay) DSOCMRDADDRVALID = DSOCMRDADDRVALID_delay;
assign #(out_delay) ISOCMBRAMEN = ISOCMBRAMEN_delay;
assign #(out_delay) ISOCMBRAMEVENWRITEEN = ISOCMBRAMEVENWRITEEN_delay;
assign #(out_delay) ISOCMBRAMODDWRITEEN = ISOCMBRAMODDWRITEEN_delay;
assign #(out_delay) ISOCMDCRBRAMEVENEN = ISOCMDCRBRAMEVENEN_delay;
assign #(out_delay) ISOCMDCRBRAMODDEN = ISOCMDCRBRAMODDEN_delay;
assign #(out_delay) ISOCMDCRBRAMRDSELECT = ISOCMDCRBRAMRDSELECT_delay;
assign #(out_delay) ISOCMBRAMRDABUS[8:28] = ISOCMBRAMRDABUS_delay[8:28];
assign #(out_delay) ISOCMBRAMWRABUS[8:28] = ISOCMBRAMWRABUS_delay[8:28];
assign #(out_delay) ISOCMBRAMWRDBUS[0:31] = ISOCMBRAMWRDBUS_delay[0:31];
assign #(out_delay) C405DBGLOADDATAONAPUDBUS = C405DBGLOADDATAONAPUDBUS_delay;
assign #(out_delay) APUFCMINSTRUCTION[0:31] = APUFCMINSTRUCTION_delay[0:31];
assign #(out_delay) APUFCMRADATA[0:31] = APUFCMRADATA_delay[0:31];
assign #(out_delay) APUFCMRBDATA[0:31] = APUFCMRBDATA_delay[0:31];
assign #(out_delay) APUFCMLOADDATA[0:31] = APUFCMLOADDATA_delay[0:31];
assign #(out_delay) APUFCMLOADBYTEEN[0:3] = APUFCMLOADBYTEEN_delay[0:3];
assign #(out_delay) APUFCMINSTRVALID = APUFCMINSTRVALID_delay;
assign #(out_delay) APUFCMOPERANDVALID = APUFCMOPERANDVALID_delay;
assign #(out_delay) APUFCMLOADDVALID = APUFCMLOADDVALID_delay;
assign #(out_delay) APUFCMFLUSH = APUFCMFLUSH_delay;
assign #(out_delay) APUFCMWRITEBACKOK = APUFCMWRITEBACKOK_delay;
assign #(out_delay) APUFCMENDIAN = APUFCMENDIAN_delay;
assign #(out_delay) APUFCMXERCA = APUFCMXERCA_delay;
assign #(out_delay) APUFCMDECODED = APUFCMDECODED_delay;
assign #(out_delay) APUFCMDECUDI[0:2] = APUFCMDECUDI_delay[0:2];
assign #(out_delay) APUFCMDECUDIVALID = APUFCMDECUDIVALID_delay;

wire	FPGA_CCLK;
wire	FPGA_BUS_RESET;
wire	FPGA_GSR;
wire	FPGA_GWE;
wire	FPGA_GHIGHB;
wire	GSR_OR;

reg	FPGA_POR;
reg	FPGA_CCLK_REG;

tri0	GSR = glbl.GSR;

`ifdef STARTUP_BLK
assign	FPGA_CCLK	= TESTBENCH.FPGA_cclk;
assign	FPGA_BUS_RESET	= TESTBENCH.FPGA_bus_reset;
assign	GSR_OR	= TESTBENCH.FPGA_gsr;
assign	FPGA_GWE	= TESTBENCH.FPGA_gwe;
assign	FPGA_GHIGHB	= TESTBENCH.FPGA_ghigh_b;
`else

FPGA_startup_VIRTEX4 start_blk(
	.bus_reset (FPGA_BUS_RESET),
	.ghigh_b (FPGA_GHIGHB),
	.gsr (FPGA_GSR),
	.done (),
	.gwe (FPGA_GWE),
	.gts_b (),
	.shutdown (1'b0),
	.cclk (FPGA_CCLK),
	.por (FPGA_POR)
);

or IGSR_OR (GSR_OR, FPGA_GSR, GSR);

`define Loc_FPGA_POR_TIME_VIRTEX4 1000 // FPGA Power-On Reset time

// Generate FPGA CCLK
always
	#5000 FPGA_CCLK_REG = ~FPGA_CCLK_REG;

assign	FPGA_CCLK = FPGA_CCLK_REG;

initial begin
	FPGA_CCLK_REG = 0;
	FPGA_POR = 1'b1;
	#(`Loc_FPGA_POR_TIME_VIRTEX4) FPGA_POR = 1'b0;
end

`endif // STARTUP_BLK

wire FPGA_BUS_RESET_delay;
wire GSR_delay;
wire FPGA_GWE_delay;
wire FPGA_GHIGHB_delay;

assign #(in_delay) FPGA_BUS_RESET_delay = FPGA_BUS_RESET;
assign #(in_delay) GSR_delay = GSR_OR;
assign #(in_delay) FPGA_GWE_delay = FPGA_GWE;
assign #(in_delay) FPGA_GHIGHB_delay = FPGA_GHIGHB;

`ifdef PROCBLK_NOSWIFT
usr_pblk_adv_cap Iusr_proc_block_cap(
`else
PPC405_ADV_SWIFT IPPC405_SWIFT(
`endif //PROCBLK_NOSWIFT

	.APUFCMDECODED (APUFCMDECODED_delay),
	.APUFCMDECUDI (APUFCMDECUDI_delay),
	.APUFCMDECUDIVALID (APUFCMDECUDIVALID_delay),
	.APUFCMENDIAN (APUFCMENDIAN_delay),
	.APUFCMFLUSH (APUFCMFLUSH_delay),
	.APUFCMINSTRUCTION (APUFCMINSTRUCTION_delay),
	.APUFCMINSTRVALID (APUFCMINSTRVALID_delay),
	.APUFCMLOADBYTEEN (APUFCMLOADBYTEEN_delay),
	.APUFCMLOADDATA (APUFCMLOADDATA_delay),
	.APUFCMLOADDVALID (APUFCMLOADDVALID_delay),
	.APUFCMOPERANDVALID (APUFCMOPERANDVALID_delay),
	.APUFCMRADATA (APUFCMRADATA_delay),
	.APUFCMRBDATA (APUFCMRBDATA_delay),
	.APUFCMWRITEBACKOK (APUFCMWRITEBACKOK_delay),
	.APUFCMXERCA (APUFCMXERCA_delay),
	.BRAMDSOCMCLK (BRAMDSOCMCLK),
	.BRAMDSOCMRDDBUS (BRAMDSOCMRDDBUS_delay),
	.BRAMISOCMCLK (BRAMISOCMCLK),
	.BRAMISOCMDCRRDDBUS (BRAMISOCMDCRRDDBUS_delay),
	.BRAMISOCMRDDBUS (BRAMISOCMRDDBUS_delay),
	.BUS_RESET (FPGA_BUS_RESET_delay),
	.C405CPMCORESLEEPREQ (C405CPMCORESLEEPREQ_delay),
	.C405CPMMSRCE (C405CPMMSRCE_delay),
	.C405CPMMSREE (C405CPMMSREE_delay),
	.C405CPMTIMERIRQ (C405CPMTIMERIRQ_delay),
	.C405CPMTIMERRESETREQ (C405CPMTIMERRESETREQ_delay),
	.C405DBGLOADDATAONAPUDBUS (C405DBGLOADDATAONAPUDBUS_delay),
	.C405DBGMSRWE (C405DBGMSRWE_delay),
	.C405DBGSTOPACK (C405DBGSTOPACK_delay),
	.C405DBGWBCOMPLETE (C405DBGWBCOMPLETE_delay),
	.C405DBGWBFULL (C405DBGWBFULL_delay),
	.C405DBGWBIAR (C405DBGWBIAR_delay),
	.C405JTGCAPTUREDR (C405JTGCAPTUREDR_delay),
	.C405JTGEXTEST (C405JTGEXTEST_delay),
	.C405JTGPGMOUT (C405JTGPGMOUT_delay),
	.C405JTGSHIFTDR (C405JTGSHIFTDR_delay),
	.C405JTGTDO (C405JTGTDO_delay),
	.C405JTGTDOEN (C405JTGTDOEN_delay),
	.C405JTGUPDATEDR (C405JTGUPDATEDR_delay),
	.C405PLBDCUABORT (C405PLBDCUABORT_delay),
	.C405PLBDCUABUS (C405PLBDCUABUS_delay),
	.C405PLBDCUBE (C405PLBDCUBE_delay),
	.C405PLBDCUCACHEABLE (C405PLBDCUCACHEABLE_delay),
	.C405PLBDCUGUARDED (C405PLBDCUGUARDED_delay),
	.C405PLBDCUPRIORITY (C405PLBDCUPRIORITY_delay),
	.C405PLBDCUREQUEST (C405PLBDCUREQUEST_delay),
	.C405PLBDCURNW (C405PLBDCURNW_delay),
	.C405PLBDCUSIZE2 (C405PLBDCUSIZE2_delay),
	.C405PLBDCUU0ATTR (C405PLBDCUU0ATTR_delay),
	.C405PLBDCUWRDBUS (C405PLBDCUWRDBUS_delay),
	.C405PLBDCUWRITETHRU (C405PLBDCUWRITETHRU_delay),
	.C405PLBICUABORT (C405PLBICUABORT_delay),
	.C405PLBICUABUS (C405PLBICUABUS_delay),
	.C405PLBICUCACHEABLE (C405PLBICUCACHEABLE_delay),
	.C405PLBICUPRIORITY (C405PLBICUPRIORITY_delay),
	.C405PLBICUREQUEST (C405PLBICUREQUEST_delay),
	.C405PLBICUSIZE (C405PLBICUSIZE_delay),
	.C405PLBICUU0ATTR (C405PLBICUU0ATTR_delay),
	.C405RSTCHIPRESETREQ (C405RSTCHIPRESETREQ_delay),
	.C405RSTCORERESETREQ (C405RSTCORERESETREQ_delay),
	.C405RSTSYSRESETREQ (C405RSTSYSRESETREQ_delay),
	.C405TRCCYCLE (C405TRCCYCLE_delay),
	.C405TRCEVENEXECUTIONSTATUS (C405TRCEVENEXECUTIONSTATUS_delay),
	.C405TRCODDEXECUTIONSTATUS (C405TRCODDEXECUTIONSTATUS_delay),
	.C405TRCTRACESTATUS (C405TRCTRACESTATUS_delay),
	.C405TRCTRIGGEREVENTOUT (C405TRCTRIGGEREVENTOUT_delay),
	.C405TRCTRIGGEREVENTTYPE (C405TRCTRIGGEREVENTTYPE_delay),
	.C405XXXMACHINECHECK (C405XXXMACHINECHECK_delay),
	.CFG_MCLK (FPGA_CCLK),
	.CPMC405CLOCK (CPMC405CLOCK),
	.CPMC405CORECLKINACTIVE (CPMC405CORECLKINACTIVE_delay),
	.CPMC405CPUCLKEN (CPMC405CPUCLKEN_delay),
	.CPMC405JTAGCLKEN (CPMC405JTAGCLKEN_delay),
	.CPMC405SYNCBYPASS (CPMC405SYNCBYPASS_delay),
	.CPMC405TIMERCLKEN (CPMC405TIMERCLKEN_delay),
	.CPMC405TIMERTICK (CPMC405TIMERTICK_delay),
	.CPMDCRCLK (CPMDCRCLK),
	.CPMFCMCLK (CPMFCMCLK),
	.DBGC405DEBUGHALT (DBGC405DEBUGHALT_delay),
	.DBGC405EXTBUSHOLDACK (DBGC405EXTBUSHOLDACK_delay),
	.DBGC405UNCONDDEBUGEVENT (DBGC405UNCONDDEBUGEVENT_delay),
	.DCREMACABUS (DCREMACABUS_delay),
	.DCREMACCLK (DCREMACCLK),
	.DCREMACDBUS (DCREMACDBUS_delay),
	.DCREMACENABLER (DCREMACENABLER_delay),
	.DCREMACREAD (DCREMACREAD_delay),
	.DCREMACWRITE (DCREMACWRITE_delay),
	.DSARCVALUE (DSARCVALUE_delay),
	.DSCNTLVALUE (DSCNTLVALUE_delay),
	.DSOCMBRAMABUS (DSOCMBRAMABUS_delay),
	.DSOCMBRAMBYTEWRITE (DSOCMBRAMBYTEWRITE_delay),
	.DSOCMBRAMEN (DSOCMBRAMEN_delay),
	.DSOCMBRAMWRDBUS (DSOCMBRAMWRDBUS_delay),
	.DSOCMBUSY (DSOCMBUSY_delay),
	.DSOCMRDADDRVALID (DSOCMRDADDRVALID_delay),
	.DSOCMRWCOMPLETE (DSOCMRWCOMPLETE_delay),
	.DSOCMWRADDRVALID (DSOCMWRADDRVALID_delay),
	.EICC405CRITINPUTIRQ (EICC405CRITINPUTIRQ_delay),
	.EICC405EXTINPUTIRQ (EICC405EXTINPUTIRQ_delay),
	.EMACDCRACK (EMACDCRACK_delay),
	.EMACDCRDBUS (EMACDCRDBUS_delay),
	.EXTDCRABUS (EXTDCRABUS_delay),
	.EXTDCRACK (EXTDCRACK_delay),
	.EXTDCRDBUSIN (EXTDCRDBUSIN_delay),
	.EXTDCRDBUSOUT (EXTDCRDBUSOUT_delay),
	.EXTDCRREAD (EXTDCRREAD_delay),
	.EXTDCRWRITE (EXTDCRWRITE_delay),
	.FCMAPUCR (FCMAPUCR_delay),
	.FCMAPUDCDCREN (FCMAPUDCDCREN_delay),
	.FCMAPUDCDFORCEALIGN (FCMAPUDCDFORCEALIGN_delay),
	.FCMAPUDCDFORCEBESTEERING (FCMAPUDCDFORCEBESTEERING_delay),
	.FCMAPUDCDFPUOP (FCMAPUDCDFPUOP_delay),
	.FCMAPUDCDGPRWRITE (FCMAPUDCDGPRWRITE_delay),
	.FCMAPUDCDLDSTBYTE (FCMAPUDCDLDSTBYTE_delay),
	.FCMAPUDCDLDSTDW (FCMAPUDCDLDSTDW_delay),
	.FCMAPUDCDLDSTHW (FCMAPUDCDLDSTHW_delay),
	.FCMAPUDCDLDSTQW (FCMAPUDCDLDSTQW_delay),
	.FCMAPUDCDLDSTWD (FCMAPUDCDLDSTWD_delay),
	.FCMAPUDCDLOAD (FCMAPUDCDLOAD_delay),
	.FCMAPUDCDPRIVOP (FCMAPUDCDPRIVOP_delay),
	.FCMAPUDCDRAEN (FCMAPUDCDRAEN_delay),
	.FCMAPUDCDRBEN (FCMAPUDCDRBEN_delay),
	.FCMAPUDCDSTORE (FCMAPUDCDSTORE_delay),
	.FCMAPUDCDTRAPBE (FCMAPUDCDTRAPBE_delay),
	.FCMAPUDCDTRAPLE (FCMAPUDCDTRAPLE_delay),
	.FCMAPUDCDUPDATE (FCMAPUDCDUPDATE_delay),
	.FCMAPUDCDXERCAEN (FCMAPUDCDXERCAEN_delay),
	.FCMAPUDCDXEROVEN (FCMAPUDCDXEROVEN_delay),
	.FCMAPUDECODEBUSY (FCMAPUDECODEBUSY_delay),
	.FCMAPUDONE (FCMAPUDONE_delay),
	.FCMAPUEXCEPTION (FCMAPUEXCEPTION_delay),
	.FCMAPUEXEBLOCKINGMCO (FCMAPUEXEBLOCKINGMCO_delay),
	.FCMAPUEXECRFIELD (FCMAPUEXECRFIELD_delay),
	.FCMAPUEXENONBLOCKINGMCO (FCMAPUEXENONBLOCKINGMCO_delay),
	.FCMAPUINSTRACK (FCMAPUINSTRACK_delay),
	.FCMAPULOADWAIT (FCMAPULOADWAIT_delay),
	.FCMAPURESULT (FCMAPURESULT_delay),
	.FCMAPURESULTVALID (FCMAPURESULTVALID_delay),
	.FCMAPUSLEEPNOTREADY (FCMAPUSLEEPNOTREADY_delay),
	.FCMAPUXERCA (FCMAPUXERCA_delay),
	.FCMAPUXEROV (FCMAPUXEROV_delay),
	.GHIGHB (FPGA_GHIGHB_delay),
	.GSR (GSR_delay),
	.GWE (FPGA_GWE_delay),
	.ISARCVALUE (ISARCVALUE_delay),
	.ISCNTLVALUE (ISCNTLVALUE_delay),
	.ISOCMBRAMEN (ISOCMBRAMEN_delay),
	.ISOCMBRAMEVENWRITEEN (ISOCMBRAMEVENWRITEEN_delay),
	.ISOCMBRAMODDWRITEEN (ISOCMBRAMODDWRITEEN_delay),
	.ISOCMBRAMRDABUS (ISOCMBRAMRDABUS_delay),
	.ISOCMBRAMWRABUS (ISOCMBRAMWRABUS_delay),
	.ISOCMBRAMWRDBUS (ISOCMBRAMWRDBUS_delay),
	.ISOCMDCRBRAMEVENEN (ISOCMDCRBRAMEVENEN_delay),
	.ISOCMDCRBRAMODDEN (ISOCMDCRBRAMODDEN_delay),
	.ISOCMDCRBRAMRDSELECT (ISOCMDCRBRAMRDSELECT_delay),
	.JTGC405BNDSCANTDO (JTGC405BNDSCANTDO_delay),
	.JTGC405TCK (JTGC405TCK),
	.JTGC405TDI (JTGC405TDI_delay),
	.JTGC405TMS (JTGC405TMS_delay),
	.JTGC405TRSTNEG (JTGC405TRSTNEG_delay),
	.MCBCPUCLKEN (MCBCPUCLKEN_delay),
	.MCBJTAGEN (MCBJTAGEN_delay),
	.MCBTIMEREN (MCBTIMEREN_delay),
	.MCPPCRST (MCPPCRST_delay),
	.PLBC405DCUADDRACK (PLBC405DCUADDRACK_delay),
	.PLBC405DCUBUSY (PLBC405DCUBUSY_delay),
	.PLBC405DCUERR (PLBC405DCUERR_delay),
	.PLBC405DCURDDACK (PLBC405DCURDDACK_delay),
	.PLBC405DCURDDBUS (PLBC405DCURDDBUS_delay),
	.PLBC405DCURDWDADDR (PLBC405DCURDWDADDR_delay),
	.PLBC405DCUSSIZE1 (PLBC405DCUSSIZE1_delay),
	.PLBC405DCUWRDACK (PLBC405DCUWRDACK_delay),
	.PLBC405ICUADDRACK (PLBC405ICUADDRACK_delay),
	.PLBC405ICUBUSY (PLBC405ICUBUSY_delay),
	.PLBC405ICUERR (PLBC405ICUERR_delay),
	.PLBC405ICURDDACK (PLBC405ICURDDACK_delay),
	.PLBC405ICURDDBUS (PLBC405ICURDDBUS_delay),
	.PLBC405ICURDWDADDR (PLBC405ICURDWDADDR_delay),
	.PLBC405ICUSSIZE1 (PLBC405ICUSSIZE1_delay),
	.PLBCLK (PLBCLK),
	.RSTC405RESETCHIP (RSTC405RESETCHIP_delay),
	.RSTC405RESETCORE (RSTC405RESETCORE_delay),
	.RSTC405RESETSYS (RSTC405RESETSYS_delay),
	.TIEAPUCONTROL (TIEAPUCONTROL_delay),
	.TIEAPUUDI1 (TIEAPUUDI1_delay),
	.TIEAPUUDI2 (TIEAPUUDI2_delay),
	.TIEAPUUDI3 (TIEAPUUDI3_delay),
	.TIEAPUUDI4 (TIEAPUUDI4_delay),
	.TIEAPUUDI5 (TIEAPUUDI5_delay),
	.TIEAPUUDI6 (TIEAPUUDI6_delay),
	.TIEAPUUDI7 (TIEAPUUDI7_delay),
	.TIEAPUUDI8 (TIEAPUUDI8_delay),
	.TIEC405DETERMINISTICMULT (TIEC405DETERMINISTICMULT_delay),
	.TIEC405DISOPERANDFWD (TIEC405DISOPERANDFWD_delay),
	.TIEC405MMUEN (TIEC405MMUEN_delay),
	.TIEDCRADDR (TIEDCRADDR_delay),
	.TIEPVRBIT10 (TIEPVRBIT10),
	.TIEPVRBIT11 (TIEPVRBIT11),
	.TIEPVRBIT28 (TIEPVRBIT28),
	.TIEPVRBIT29 (TIEPVRBIT29),
	.TIEPVRBIT30 (TIEPVRBIT30),
	.TIEPVRBIT31 (TIEPVRBIT31),
	.TIEPVRBIT8 (TIEPVRBIT8),
	.TIEPVRBIT9 (TIEPVRBIT9),
	.TRCC405TRACEDISABLE (TRCC405TRACEDISABLE_delay),
	.TRCC405TRIGGEREVENTIN (TRCC405TRIGGEREVENTIN_delay)
);

endmodule

module FPGA_startup_VIRTEX4 (bus_reset, ghigh_b, gsr, done, gwe, gts_b, shutdown, cclk, por);

output bus_reset;
output ghigh_b;
output gsr;
output done;
output gwe;
output gts_b;

input shutdown;
input cclk, por;

reg bus_reset, abus_reset;
reg ghigh_b, aghigh_b;
reg gsr, agsr;
reg done, adone;
reg gwe, agwe;
reg gts_b, agts_b;

reg [7:0] count;

always @ (posedge cclk or posedge por) begin
	if (por) count <= {8{1'b0}};
	else if (shutdown &&(count > {8{1'b0}})) count = count - 1;
	else if (!shutdown &&(count < {8'hFF})) count = count + 1;
end

always @ (posedge cclk or posedge por) begin
	if (por) begin
		{bus_reset,ghigh_b,gsr,done,gwe,gts_b} <= 6'b100000;
	end
	else begin
		{bus_reset,ghigh_b,gsr,done,gwe,gts_b} <= {abus_reset,aghigh_b,agsr,adone,agwe,agts_b};
	end
end

always @ (count) begin
	// defaults

	abus_reset = 1;
	aghigh_b = 0;
	agsr = 0;
	adone = 0;
	agwe = 0;
	agts_b = 0;

	// Trip times are in order for default sequence.
	if (count >= 8'h02) abus_reset = 0;
	if (count == 8'h17 || count == 8'h18) agsr = 1;
	if (count > 8'h27) aghigh_b = 1;
	if (count > 8'h31) adone = 1;
	if (count == 8'h33 || count == 8'h34) agsr = 1;
	if (count > 8'h36) agwe = 1;
	if (count > 8'h37) agts_b = 1;
end

endmodule // FPGA_startup
