// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/USR_ACCESS_VIRTEX4.v,v 1.1.4.4 2004/05/12 19:07:23 patrickp Exp $

`timescale  100 ps / 10 ps

module USR_ACCESS_VIRTEX4 (DATA, DATAVALID);

    output [31:0] DATA;
    output DATAVALID;

endmodule // USR_ACCESS_VIRTEX4
