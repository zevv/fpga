// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/TIMEGRP.v,v 1.8.22.1 2003/11/18 20:41:40 wloo Exp $

/*

FUNCTION	: TIMEGRP dummy simulation module

*/

`timescale  100 ps / 10 ps


module TIMEGRP ();

endmodule

