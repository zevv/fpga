// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/TIMESPEC.v,v 1.8.22.1 2003/11/18 20:41:40 wloo Exp $

/*

FUNCTION	: TIMESPEC dummy simulation module

*/

`timescale  100 ps / 10 ps


module TIMESPEC ();

endmodule

