// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/CONFIG.v,v 1.8.22.1 2003/11/18 20:41:33 wloo Exp $

/*

FUNCTION	: CONFIG dummy simulation module

*/

`timescale  100 ps / 10 ps


module CONFIG ();

endmodule

