// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/EMAC.v,v 1.1.4.6 2004/09/15 15:59:30 patrickp Exp $

`timescale 1 ps / 1 ps 

module EMAC (
	DCRHOSTDONEIR,
	EMAC0CLIENTANINTERRUPT,
	EMAC0CLIENTRXBADFRAME,
	EMAC0CLIENTRXCLIENTCLKOUT,
	EMAC0CLIENTRXD,
	EMAC0CLIENTRXDVLD,
	EMAC0CLIENTRXDVLDMSW,
	EMAC0CLIENTRXDVREG6,
	EMAC0CLIENTRXFRAMEDROP,
	EMAC0CLIENTRXGOODFRAME,
	EMAC0CLIENTRXSTATS,
	EMAC0CLIENTRXSTATSBYTEVLD,
	EMAC0CLIENTRXSTATSVLD,
	EMAC0CLIENTTXACK,
	EMAC0CLIENTTXCLIENTCLKOUT,
	EMAC0CLIENTTXCOLLISION,
	EMAC0CLIENTTXGMIIMIICLKOUT,
	EMAC0CLIENTTXRETRANSMIT,
	EMAC0CLIENTTXSTATS,
	EMAC0CLIENTTXSTATSBYTEVLD,
	EMAC0CLIENTTXSTATSVLD,
	EMAC0PHYENCOMMAALIGN,
	EMAC0PHYLOOPBACKMSB,
	EMAC0PHYMCLKOUT,
	EMAC0PHYMDOUT,
	EMAC0PHYMDTRI,
	EMAC0PHYMGTRXRESET,
	EMAC0PHYMGTTXRESET,
	EMAC0PHYPOWERDOWN,
	EMAC0PHYSYNCACQSTATUS,
	EMAC0PHYTXCHARDISPMODE,
	EMAC0PHYTXCHARDISPVAL,
	EMAC0PHYTXCHARISK,
	EMAC0PHYTXCLK,
	EMAC0PHYTXD,
	EMAC0PHYTXEN,
	EMAC0PHYTXER,
	EMAC1CLIENTANINTERRUPT,
	EMAC1CLIENTRXBADFRAME,
	EMAC1CLIENTRXCLIENTCLKOUT,
	EMAC1CLIENTRXD,
	EMAC1CLIENTRXDVLD,
	EMAC1CLIENTRXDVLDMSW,
	EMAC1CLIENTRXDVREG6,
	EMAC1CLIENTRXFRAMEDROP,
	EMAC1CLIENTRXGOODFRAME,
	EMAC1CLIENTRXSTATS,
	EMAC1CLIENTRXSTATSBYTEVLD,
	EMAC1CLIENTRXSTATSVLD,
	EMAC1CLIENTTXACK,
	EMAC1CLIENTTXCLIENTCLKOUT,
	EMAC1CLIENTTXCOLLISION,
	EMAC1CLIENTTXGMIIMIICLKOUT,
	EMAC1CLIENTTXRETRANSMIT,
	EMAC1CLIENTTXSTATS,
	EMAC1CLIENTTXSTATSBYTEVLD,
	EMAC1CLIENTTXSTATSVLD,
	EMAC1PHYENCOMMAALIGN,
	EMAC1PHYLOOPBACKMSB,
	EMAC1PHYMCLKOUT,
	EMAC1PHYMDOUT,
	EMAC1PHYMDTRI,
	EMAC1PHYMGTRXRESET,
	EMAC1PHYMGTTXRESET,
	EMAC1PHYPOWERDOWN,
	EMAC1PHYSYNCACQSTATUS,
	EMAC1PHYTXCHARDISPMODE,
	EMAC1PHYTXCHARDISPVAL,
	EMAC1PHYTXCHARISK,
	EMAC1PHYTXCLK,
	EMAC1PHYTXD,
	EMAC1PHYTXEN,
	EMAC1PHYTXER,
	EMACDCRACK,
	EMACDCRDBUS,
	HOSTMIIMRDY,
	HOSTRDDATA,
	CLIENTEMAC0DCMLOCKED,
	CLIENTEMAC0PAUSEREQ,
	CLIENTEMAC0PAUSEVAL,
	CLIENTEMAC0RXCLIENTCLKIN,
	CLIENTEMAC0TXCLIENTCLKIN,
	CLIENTEMAC0TXD,
	CLIENTEMAC0TXDVLD,
	CLIENTEMAC0TXDVLDMSW,
	CLIENTEMAC0TXFIRSTBYTE,
	CLIENTEMAC0TXGMIIMIICLKIN,
	CLIENTEMAC0TXIFGDELAY,
	CLIENTEMAC0TXUNDERRUN,
	CLIENTEMAC1DCMLOCKED,
	CLIENTEMAC1PAUSEREQ,
	CLIENTEMAC1PAUSEVAL,
	CLIENTEMAC1RXCLIENTCLKIN,
	CLIENTEMAC1TXCLIENTCLKIN,
	CLIENTEMAC1TXD,
	CLIENTEMAC1TXDVLD,
	CLIENTEMAC1TXDVLDMSW,
	CLIENTEMAC1TXFIRSTBYTE,
	CLIENTEMAC1TXGMIIMIICLKIN,
	CLIENTEMAC1TXIFGDELAY,
	CLIENTEMAC1TXUNDERRUN,
	DCREMACABUS,
	DCREMACCLK,
	DCREMACDBUS,
	DCREMACENABLE,
	DCREMACREAD,
	DCREMACWRITE,
	HOSTADDR,
	HOSTCLK,
	HOSTEMAC1SEL,
	HOSTMIIMSEL,
	HOSTOPCODE,
	HOSTREQ,
	HOSTWRDATA,
	PHYEMAC0COL,
	PHYEMAC0CRS,
	PHYEMAC0GTXCLK,
	PHYEMAC0MCLKIN,
	PHYEMAC0MDIN,
	PHYEMAC0MIITXCLK,
	PHYEMAC0PHYAD,
	PHYEMAC0RXBUFERR,
	PHYEMAC0RXBUFSTATUS,
	PHYEMAC0RXCHARISCOMMA,
	PHYEMAC0RXCHARISK,
	PHYEMAC0RXCHECKINGCRC,
	PHYEMAC0RXCLK,
	PHYEMAC0RXCLKCORCNT,
	PHYEMAC0RXCOMMADET,
	PHYEMAC0RXD,
	PHYEMAC0RXDISPERR,
	PHYEMAC0RXDV,
	PHYEMAC0RXER,
	PHYEMAC0RXLOSSOFSYNC,
	PHYEMAC0RXNOTINTABLE,
	PHYEMAC0RXRUNDISP,
	PHYEMAC0SIGNALDET,
	PHYEMAC0TXBUFERR,
	PHYEMAC1COL,
	PHYEMAC1CRS,
	PHYEMAC1GTXCLK,
	PHYEMAC1MCLKIN,
	PHYEMAC1MDIN,
	PHYEMAC1MIITXCLK,
	PHYEMAC1PHYAD,
	PHYEMAC1RXBUFERR,
	PHYEMAC1RXBUFSTATUS,
	PHYEMAC1RXCHARISCOMMA,
	PHYEMAC1RXCHARISK,
	PHYEMAC1RXCHECKINGCRC,
	PHYEMAC1RXCLK,
	PHYEMAC1RXCLKCORCNT,
	PHYEMAC1RXCOMMADET,
	PHYEMAC1RXD,
	PHYEMAC1RXDISPERR,
	PHYEMAC1RXDV,
	PHYEMAC1RXER,
	PHYEMAC1RXLOSSOFSYNC,
	PHYEMAC1RXNOTINTABLE,
	PHYEMAC1RXRUNDISP,
	PHYEMAC1SIGNALDET,
	PHYEMAC1TXBUFERR,
	RESET,
	TIEEMAC0CONFIGVEC,
	TIEEMAC0UNICASTADDR,
	TIEEMAC1CONFIGVEC,
	TIEEMAC1UNICASTADDR
);

parameter in_delay = 100;
parameter out_delay = 100;

output DCRHOSTDONEIR;
output EMAC0CLIENTANINTERRUPT;
output EMAC0CLIENTRXBADFRAME;
output EMAC0CLIENTRXCLIENTCLKOUT;
output EMAC0CLIENTRXDVLD;
output EMAC0CLIENTRXDVLDMSW;
output EMAC0CLIENTRXDVREG6;
output EMAC0CLIENTRXFRAMEDROP;
output EMAC0CLIENTRXGOODFRAME;
output EMAC0CLIENTRXSTATSBYTEVLD;
output EMAC0CLIENTRXSTATSVLD;
output EMAC0CLIENTTXACK;
output EMAC0CLIENTTXCLIENTCLKOUT;
output EMAC0CLIENTTXCOLLISION;
output EMAC0CLIENTTXGMIIMIICLKOUT;
output EMAC0CLIENTTXRETRANSMIT;
output EMAC0CLIENTTXSTATS;
output EMAC0CLIENTTXSTATSBYTEVLD;
output EMAC0CLIENTTXSTATSVLD;
output EMAC0PHYENCOMMAALIGN;
output EMAC0PHYLOOPBACKMSB;
output EMAC0PHYMCLKOUT;
output EMAC0PHYMDOUT;
output EMAC0PHYMDTRI;
output EMAC0PHYMGTRXRESET;
output EMAC0PHYMGTTXRESET;
output EMAC0PHYPOWERDOWN;
output EMAC0PHYSYNCACQSTATUS;
output EMAC0PHYTXCHARDISPMODE;
output EMAC0PHYTXCHARDISPVAL;
output EMAC0PHYTXCHARISK;
output EMAC0PHYTXCLK;
output EMAC0PHYTXEN;
output EMAC0PHYTXER;
output EMAC1CLIENTANINTERRUPT;
output EMAC1CLIENTRXBADFRAME;
output EMAC1CLIENTRXCLIENTCLKOUT;
output EMAC1CLIENTRXDVLD;
output EMAC1CLIENTRXDVLDMSW;
output EMAC1CLIENTRXDVREG6;
output EMAC1CLIENTRXFRAMEDROP;
output EMAC1CLIENTRXGOODFRAME;
output EMAC1CLIENTRXSTATSBYTEVLD;
output EMAC1CLIENTRXSTATSVLD;
output EMAC1CLIENTTXACK;
output EMAC1CLIENTTXCLIENTCLKOUT;
output EMAC1CLIENTTXCOLLISION;
output EMAC1CLIENTTXGMIIMIICLKOUT;
output EMAC1CLIENTTXRETRANSMIT;
output EMAC1CLIENTTXSTATS;
output EMAC1CLIENTTXSTATSBYTEVLD;
output EMAC1CLIENTTXSTATSVLD;
output EMAC1PHYENCOMMAALIGN;
output EMAC1PHYLOOPBACKMSB;
output EMAC1PHYMCLKOUT;
output EMAC1PHYMDOUT;
output EMAC1PHYMDTRI;
output EMAC1PHYMGTRXRESET;
output EMAC1PHYMGTTXRESET;
output EMAC1PHYPOWERDOWN;
output EMAC1PHYSYNCACQSTATUS;
output EMAC1PHYTXCHARDISPMODE;
output EMAC1PHYTXCHARDISPVAL;
output EMAC1PHYTXCHARISK;
output EMAC1PHYTXCLK;
output EMAC1PHYTXEN;
output EMAC1PHYTXER;
output EMACDCRACK;
output HOSTMIIMRDY;
output [0:31] EMACDCRDBUS;
output [15:0] EMAC0CLIENTRXD;
output [15:0] EMAC1CLIENTRXD;
output [31:0] HOSTRDDATA;
output [6:0] EMAC0CLIENTRXSTATS;
output [6:0] EMAC1CLIENTRXSTATS;
output [7:0] EMAC0PHYTXD;
output [7:0] EMAC1PHYTXD;

input CLIENTEMAC0DCMLOCKED;
input CLIENTEMAC0PAUSEREQ;
input CLIENTEMAC0RXCLIENTCLKIN;
input CLIENTEMAC0TXCLIENTCLKIN;
input CLIENTEMAC0TXDVLD;
input CLIENTEMAC0TXDVLDMSW;
input CLIENTEMAC0TXFIRSTBYTE;
input CLIENTEMAC0TXGMIIMIICLKIN;
input CLIENTEMAC0TXUNDERRUN;
input CLIENTEMAC1DCMLOCKED;
input CLIENTEMAC1PAUSEREQ;
input CLIENTEMAC1RXCLIENTCLKIN;
input CLIENTEMAC1TXCLIENTCLKIN;
input CLIENTEMAC1TXDVLD;
input CLIENTEMAC1TXDVLDMSW;
input CLIENTEMAC1TXFIRSTBYTE;
input CLIENTEMAC1TXGMIIMIICLKIN;
input CLIENTEMAC1TXUNDERRUN;
input DCREMACCLK;
input DCREMACENABLE;
input DCREMACREAD;
input DCREMACWRITE;
input HOSTCLK;
input HOSTEMAC1SEL;
input HOSTMIIMSEL;
input HOSTREQ;
input PHYEMAC0COL;
input PHYEMAC0CRS;
input PHYEMAC0GTXCLK;
input PHYEMAC0MCLKIN;
input PHYEMAC0MDIN;
input PHYEMAC0MIITXCLK;
input PHYEMAC0RXBUFERR;
input PHYEMAC0RXCHARISCOMMA;
input PHYEMAC0RXCHARISK;
input PHYEMAC0RXCHECKINGCRC;
input PHYEMAC0RXCLK;
input PHYEMAC0RXCOMMADET;
input PHYEMAC0RXDISPERR;
input PHYEMAC0RXDV;
input PHYEMAC0RXER;
input PHYEMAC0RXNOTINTABLE;
input PHYEMAC0RXRUNDISP;
input PHYEMAC0SIGNALDET;
input PHYEMAC0TXBUFERR;
input PHYEMAC1COL;
input PHYEMAC1CRS;
input PHYEMAC1GTXCLK;
input PHYEMAC1MCLKIN;
input PHYEMAC1MDIN;
input PHYEMAC1MIITXCLK;
input PHYEMAC1RXBUFERR;
input PHYEMAC1RXCHARISCOMMA;
input PHYEMAC1RXCHARISK;
input PHYEMAC1RXCHECKINGCRC;
input PHYEMAC1RXCLK;
input PHYEMAC1RXCOMMADET;
input PHYEMAC1RXDISPERR;
input PHYEMAC1RXDV;
input PHYEMAC1RXER;
input PHYEMAC1RXNOTINTABLE;
input PHYEMAC1RXRUNDISP;
input PHYEMAC1SIGNALDET;
input PHYEMAC1TXBUFERR;
input RESET;
input [0:31] DCREMACDBUS;
input [15:0] CLIENTEMAC0PAUSEVAL;
input [15:0] CLIENTEMAC0TXD;
input [15:0] CLIENTEMAC1PAUSEVAL;
input [15:0] CLIENTEMAC1TXD;
input [1:0] HOSTOPCODE;
input [1:0] PHYEMAC0RXBUFSTATUS;
input [1:0] PHYEMAC0RXLOSSOFSYNC;
input [1:0] PHYEMAC1RXBUFSTATUS;
input [1:0] PHYEMAC1RXLOSSOFSYNC;
input [2:0] PHYEMAC0RXCLKCORCNT;
input [2:0] PHYEMAC1RXCLKCORCNT;
input [31:0] HOSTWRDATA;
input [47:0] TIEEMAC0UNICASTADDR;
input [47:0] TIEEMAC1UNICASTADDR;
input [4:0] PHYEMAC0PHYAD;
input [4:0] PHYEMAC1PHYAD;
input [79:0] TIEEMAC0CONFIGVEC;
input [79:0] TIEEMAC1CONFIGVEC;
input [7:0] CLIENTEMAC0TXIFGDELAY;
input [7:0] CLIENTEMAC1TXIFGDELAY;
input [7:0] PHYEMAC0RXD;
input [7:0] PHYEMAC1RXD;
input [8:9] DCREMACABUS;
input [9:0] HOSTADDR;

wire CLIENTEMAC0DCMLOCKED_delay; 
wire CLIENTEMAC0PAUSEREQ_delay;
wire CLIENTEMAC0TXDVLDMSW_delay;
wire CLIENTEMAC0TXDVLD_delay;
wire CLIENTEMAC0TXFIRSTBYTE_delay;
wire CLIENTEMAC0TXUNDERRUN_delay;
wire CLIENTEMAC1DCMLOCKED_delay; 
wire CLIENTEMAC1PAUSEREQ_delay;
wire CLIENTEMAC1TXDVLDMSW_delay;
wire CLIENTEMAC1TXDVLD_delay;
wire CLIENTEMAC1TXFIRSTBYTE_delay;
wire CLIENTEMAC1TXUNDERRUN_delay;
wire DCREMACENABLE_delay; // HOSTUSEDCR;
wire DCREMACREAD_delay;
wire DCREMACWRITE_delay;
wire DCRHOSTDONEIR; 
wire DCRHOSTDONEIR_delay; 
wire EMAC0CLIENTANINTERRUPT; 
wire EMAC0CLIENTANINTERRUPT_delay; 
wire EMAC0CLIENTRXBADFRAME;
wire EMAC0CLIENTRXBADFRAME_delay;
wire EMAC0CLIENTRXCLIENTCLKOUT; 
wire EMAC0CLIENTRXDVLD;
wire EMAC0CLIENTRXDVLDMSW;
wire EMAC0CLIENTRXDVLDMSW_delay;
wire EMAC0CLIENTRXDVLD_delay;
wire EMAC0CLIENTRXDVREG6;
wire EMAC0CLIENTRXDVREG6_delay;
wire EMAC0CLIENTRXFRAMEDROP;
wire EMAC0CLIENTRXFRAMEDROP_delay;
wire EMAC0CLIENTRXGOODFRAME;
wire EMAC0CLIENTRXGOODFRAME_delay;
wire EMAC0CLIENTRXSTATSBYTEVLD;
wire EMAC0CLIENTRXSTATSBYTEVLD_delay;
wire EMAC0CLIENTRXSTATSVLD;
wire EMAC0CLIENTRXSTATSVLD_delay;
wire EMAC0CLIENTTXACK;
wire EMAC0CLIENTTXACK_delay;
wire EMAC0CLIENTTXCLIENTCLKOUT; 
wire EMAC0CLIENTTXCOLLISION;
wire EMAC0CLIENTTXCOLLISION_delay;
wire EMAC0CLIENTTXGMIIMIICLKOUT; 
wire EMAC0CLIENTTXRETRANSMIT;
wire EMAC0CLIENTTXRETRANSMIT_delay;
wire EMAC0CLIENTTXSTATS;
wire EMAC0CLIENTTXSTATSBYTEVLD;
wire EMAC0CLIENTTXSTATSBYTEVLD_delay;
wire EMAC0CLIENTTXSTATSVLD;
wire EMAC0CLIENTTXSTATSVLD_delay;
wire EMAC0CLIENTTXSTATS_delay;
wire EMAC0PHYENCOMMAALIGN; 
wire EMAC0PHYENCOMMAALIGN_delay; 
wire EMAC0PHYLOOPBACKMSB;
wire EMAC0PHYLOOPBACKMSB_delay;
wire EMAC0PHYMCLKOUT;
wire EMAC0PHYMCLKOUT_delay;
wire EMAC0PHYMDOUT;
wire EMAC0PHYMDOUT_delay;
wire EMAC0PHYMDTRI;
wire EMAC0PHYMDTRI_delay;
wire EMAC0PHYMGTRXRESET; 
wire EMAC0PHYMGTRXRESET_delay; 
wire EMAC0PHYMGTTXRESET; 
wire EMAC0PHYMGTTXRESET_delay; 
wire EMAC0PHYPOWERDOWN; 
wire EMAC0PHYPOWERDOWN_delay; 
wire EMAC0PHYSYNCACQSTATUS; 
wire EMAC0PHYSYNCACQSTATUS_delay; 
wire EMAC0PHYTXCHARDISPMODE;
wire EMAC0PHYTXCHARDISPMODE_delay;
wire EMAC0PHYTXCHARDISPVAL;
wire EMAC0PHYTXCHARDISPVAL_delay;
wire EMAC0PHYTXCHARISK;
wire EMAC0PHYTXCHARISK_delay;
wire EMAC0PHYTXCLK; 
wire EMAC0PHYTXEN;
wire EMAC0PHYTXEN_delay;
wire EMAC0PHYTXER;
wire EMAC0PHYTXER_delay;
wire EMAC1CLIENTANINTERRUPT; 
wire EMAC1CLIENTANINTERRUPT_delay; 
wire EMAC1CLIENTRXBADFRAME;
wire EMAC1CLIENTRXBADFRAME_delay;
wire EMAC1CLIENTRXCLIENTCLKOUT; 
wire EMAC1CLIENTRXDVLD;
wire EMAC1CLIENTRXDVLDMSW;
wire EMAC1CLIENTRXDVLDMSW_delay;
wire EMAC1CLIENTRXDVLD_delay;
wire EMAC1CLIENTRXDVREG6;
wire EMAC1CLIENTRXDVREG6_delay;
wire EMAC1CLIENTRXFRAMEDROP;
wire EMAC1CLIENTRXFRAMEDROP_delay;
wire EMAC1CLIENTRXGOODFRAME;
wire EMAC1CLIENTRXGOODFRAME_delay;
wire EMAC1CLIENTRXSTATSBYTEVLD;
wire EMAC1CLIENTRXSTATSBYTEVLD_delay;
wire EMAC1CLIENTRXSTATSVLD;
wire EMAC1CLIENTRXSTATSVLD_delay;
wire EMAC1CLIENTTXACK;
wire EMAC1CLIENTTXACK_delay;
wire EMAC1CLIENTTXCLIENTCLKOUT; 
wire EMAC1CLIENTTXCOLLISION;
wire EMAC1CLIENTTXCOLLISION_delay;
wire EMAC1CLIENTTXGMIIMIICLKOUT; 
wire EMAC1CLIENTTXRETRANSMIT;
wire EMAC1CLIENTTXRETRANSMIT_delay;
wire EMAC1CLIENTTXSTATS;
wire EMAC1CLIENTTXSTATSBYTEVLD;
wire EMAC1CLIENTTXSTATSBYTEVLD_delay;
wire EMAC1CLIENTTXSTATSVLD;
wire EMAC1CLIENTTXSTATSVLD_delay;
wire EMAC1CLIENTTXSTATS_delay;
wire EMAC1PHYENCOMMAALIGN; 
wire EMAC1PHYENCOMMAALIGN_delay; 
wire EMAC1PHYLOOPBACKMSB;
wire EMAC1PHYLOOPBACKMSB_delay;
wire EMAC1PHYMCLKOUT;
wire EMAC1PHYMCLKOUT_delay;
wire EMAC1PHYMDOUT;
wire EMAC1PHYMDOUT_delay;
wire EMAC1PHYMDTRI;
wire EMAC1PHYMDTRI_delay;
wire EMAC1PHYMGTRXRESET; 
wire EMAC1PHYMGTRXRESET_delay; 
wire EMAC1PHYMGTTXRESET; 
wire EMAC1PHYMGTTXRESET_delay; 
wire EMAC1PHYPOWERDOWN; 
wire EMAC1PHYPOWERDOWN_delay; 
wire EMAC1PHYSYNCACQSTATUS; 
wire EMAC1PHYSYNCACQSTATUS_delay; 
wire EMAC1PHYTXCHARDISPMODE;
wire EMAC1PHYTXCHARDISPMODE_delay;
wire EMAC1PHYTXCHARDISPVAL;
wire EMAC1PHYTXCHARDISPVAL_delay;
wire EMAC1PHYTXCHARISK;
wire EMAC1PHYTXCHARISK_delay;
wire EMAC1PHYTXCLK;
wire EMAC1PHYTXEN;
wire EMAC1PHYTXEN_delay;
wire EMAC1PHYTXER;
wire EMAC1PHYTXER_delay;
wire EMACDCRACK;
wire EMACDCRACK_delay;
wire HOSTEMAC1SEL_delay;
wire HOSTMIIMRDY;
wire HOSTMIIMRDY_delay;
wire HOSTMIIMSEL_delay;
wire HOSTREQ_delay;
wire PHYEMAC0COL_delay;
wire PHYEMAC0CRS_delay;
wire PHYEMAC0MCLKIN_delay;
wire PHYEMAC0MDIN_delay;
wire PHYEMAC0RXBUFERR_delay;
wire PHYEMAC0RXCHARISCOMMA_delay;
wire PHYEMAC0RXCHARISK_delay;
wire PHYEMAC0RXCHECKINGCRC_delay;
wire PHYEMAC0RXCOMMADET_delay; 
wire PHYEMAC0RXDISPERR_delay;
wire PHYEMAC0RXDV_delay;
wire PHYEMAC0RXER_delay;
wire PHYEMAC0RXNOTINTABLE_delay;
wire PHYEMAC0RXRUNDISP_delay;
wire PHYEMAC0SIGNALDET_delay; 
wire PHYEMAC0TXBUFERR_delay;
wire PHYEMAC1COL_delay;
wire PHYEMAC1CRS_delay;
wire PHYEMAC1MCLKIN_delay;
wire PHYEMAC1MDIN_delay;
wire PHYEMAC1RXBUFERR_delay;
wire PHYEMAC1RXCHARISCOMMA_delay;
wire PHYEMAC1RXCHARISK_delay;
wire PHYEMAC1RXCHECKINGCRC_delay;
wire PHYEMAC1RXCOMMADET_delay; 
wire PHYEMAC1RXDISPERR_delay;
wire PHYEMAC1RXDV_delay;
wire PHYEMAC1RXER_delay;
wire PHYEMAC1RXNOTINTABLE_delay;
wire PHYEMAC1RXRUNDISP_delay;
wire PHYEMAC1SIGNALDET_delay; 
wire PHYEMAC1TXBUFERR_delay;
wire RESET_delay;
wire [0:31] DCREMACDBUS_delay;
wire [0:31] EMACDCRDBUS;
wire [0:31] EMACDCRDBUS_delay;
wire [15:0] CLIENTEMAC0PAUSEVAL_delay;
wire [15:0] CLIENTEMAC0TXD_delay;
wire [15:0] CLIENTEMAC1PAUSEVAL_delay;
wire [15:0] CLIENTEMAC1TXD_delay;
wire [15:0] EMAC0CLIENTRXD;
wire [15:0] EMAC0CLIENTRXD_delay;
wire [15:0] EMAC1CLIENTRXD;
wire [15:0] EMAC1CLIENTRXD_delay;
wire [1:0] HOSTOPCODE_delay;
wire [1:0] PHYEMAC0RXBUFSTATUS_delay;
wire [1:0] PHYEMAC0RXLOSSOFSYNC_delay;
wire [1:0] PHYEMAC1RXBUFSTATUS_delay;
wire [1:0] PHYEMAC1RXLOSSOFSYNC_delay;
wire [2:0] PHYEMAC0RXCLKCORCNT_delay; 
wire [2:0] PHYEMAC1RXCLKCORCNT_delay; 
wire [31:0] HOSTRDDATA;
wire [31:0] HOSTRDDATA_delay;
wire [31:0] HOSTWRDATA_delay;
wire [47:0] TIEEMAC0UNICASTADDR_delay;
wire [47:0] TIEEMAC1UNICASTADDR_delay;
wire [4:0] PHYEMAC0PHYAD_delay; 
wire [4:0] PHYEMAC1PHYAD_delay;
wire [6:0] EMAC0CLIENTRXSTATS;
wire [6:0] EMAC0CLIENTRXSTATS_delay;
wire [6:0] EMAC1CLIENTRXSTATS;
wire [6:0] EMAC1CLIENTRXSTATS_delay;
wire [79:0] TIEEMAC0CONFIGVEC_delay;
wire [79:0] TIEEMAC1CONFIGVEC_delay;
wire [7:0] CLIENTEMAC0TXIFGDELAY_delay;
wire [7:0] CLIENTEMAC1TXIFGDELAY_delay;
wire [7:0] EMAC0PHYTXD;
wire [7:0] EMAC0PHYTXD_delay;
wire [7:0] EMAC1PHYTXD;
wire [7:0] EMAC1PHYTXD_delay;
wire [7:0] PHYEMAC0RXD_delay;
wire [7:0] PHYEMAC1RXD_delay;
wire [8:9] DCREMACABUS_delay; 
wire [9:0] HOSTADDR_delay;



assign #(in_delay) CLIENTEMAC0DCMLOCKED_delay = CLIENTEMAC0DCMLOCKED;
assign #(in_delay) CLIENTEMAC0PAUSEREQ_delay = CLIENTEMAC0PAUSEREQ;
assign #(in_delay) CLIENTEMAC0PAUSEVAL_delay[15:0] = CLIENTEMAC0PAUSEVAL[15:0];
assign #(in_delay) CLIENTEMAC0TXDVLDMSW_delay = CLIENTEMAC0TXDVLDMSW;
assign #(in_delay) CLIENTEMAC0TXDVLD_delay = CLIENTEMAC0TXDVLD;
assign #(in_delay) CLIENTEMAC0TXD_delay[15:0] = CLIENTEMAC0TXD[15:0];
assign #(in_delay) CLIENTEMAC0TXFIRSTBYTE_delay = CLIENTEMAC0TXFIRSTBYTE;
assign #(in_delay) CLIENTEMAC0TXIFGDELAY_delay[7:0] = CLIENTEMAC0TXIFGDELAY[7:0];
assign #(in_delay) CLIENTEMAC0TXUNDERRUN_delay = CLIENTEMAC0TXUNDERRUN;
assign #(in_delay) CLIENTEMAC1DCMLOCKED_delay = CLIENTEMAC1DCMLOCKED;
assign #(in_delay) CLIENTEMAC1PAUSEREQ_delay = CLIENTEMAC1PAUSEREQ;
assign #(in_delay) CLIENTEMAC1PAUSEVAL_delay[15:0] = CLIENTEMAC1PAUSEVAL[15:0];
assign #(in_delay) CLIENTEMAC1TXDVLDMSW_delay = CLIENTEMAC1TXDVLDMSW;
assign #(in_delay) CLIENTEMAC1TXDVLD_delay = CLIENTEMAC1TXDVLD;
assign #(in_delay) CLIENTEMAC1TXD_delay[15:0] = CLIENTEMAC1TXD[15:0];
assign #(in_delay) CLIENTEMAC1TXFIRSTBYTE_delay = CLIENTEMAC1TXFIRSTBYTE;
assign #(in_delay) CLIENTEMAC1TXIFGDELAY_delay[7:0] = CLIENTEMAC1TXIFGDELAY[7:0];
assign #(in_delay) CLIENTEMAC1TXUNDERRUN_delay = CLIENTEMAC1TXUNDERRUN;
assign #(in_delay) DCREMACABUS_delay[8:9] = DCREMACABUS[8:9];
assign #(in_delay) DCREMACDBUS_delay[0:31] = DCREMACDBUS[0:31];
assign #(in_delay) DCREMACENABLE_delay = DCREMACENABLE;
assign #(in_delay) DCREMACREAD_delay = DCREMACREAD;
assign #(in_delay) DCREMACWRITE_delay = DCREMACWRITE;
assign #(in_delay) HOSTADDR_delay[9:0] = HOSTADDR[9:0];
assign #(in_delay) HOSTEMAC1SEL_delay = HOSTEMAC1SEL;
assign #(in_delay) HOSTMIIMSEL_delay = HOSTMIIMSEL;
assign #(in_delay) HOSTOPCODE_delay[1:0] = HOSTOPCODE[1:0];
assign #(in_delay) HOSTREQ_delay = HOSTREQ;
assign #(in_delay) HOSTWRDATA_delay[31:0] = HOSTWRDATA[31:0];
assign #(in_delay) PHYEMAC0COL_delay = PHYEMAC0COL;
assign #(in_delay) PHYEMAC0CRS_delay = PHYEMAC0CRS;
assign #(in_delay) PHYEMAC0MCLKIN_delay = PHYEMAC0MCLKIN;
assign #(in_delay) PHYEMAC0MDIN_delay = PHYEMAC0MDIN;
assign #(in_delay) PHYEMAC0PHYAD_delay[4:0] = PHYEMAC0PHYAD[4:0];
assign #(in_delay) PHYEMAC0RXBUFERR_delay = PHYEMAC0RXBUFERR;
assign #(in_delay) PHYEMAC0RXBUFSTATUS_delay[1:0] = PHYEMAC0RXBUFSTATUS[1:0];
assign #(in_delay) PHYEMAC0RXCHARISCOMMA_delay = PHYEMAC0RXCHARISCOMMA;
assign #(in_delay) PHYEMAC0RXCHARISK_delay = PHYEMAC0RXCHARISK;
assign #(in_delay) PHYEMAC0RXCHECKINGCRC_delay = PHYEMAC0RXCHECKINGCRC;
assign #(in_delay) PHYEMAC0RXCLKCORCNT_delay[2:0] = PHYEMAC0RXCLKCORCNT[2:0];
assign #(in_delay) PHYEMAC0RXCOMMADET_delay = PHYEMAC0RXCOMMADET;
assign #(in_delay) PHYEMAC0RXDISPERR_delay = PHYEMAC0RXDISPERR;
assign #(in_delay) PHYEMAC0RXDV_delay = PHYEMAC0RXDV;
assign #(in_delay) PHYEMAC0RXD_delay[7:0] = PHYEMAC0RXD[7:0];
assign #(in_delay) PHYEMAC0RXER_delay = PHYEMAC0RXER;
assign #(in_delay) PHYEMAC0RXLOSSOFSYNC_delay[1:0] = PHYEMAC0RXLOSSOFSYNC[1:0];
assign #(in_delay) PHYEMAC0RXNOTINTABLE_delay = PHYEMAC0RXNOTINTABLE;
assign #(in_delay) PHYEMAC0RXRUNDISP_delay = PHYEMAC0RXRUNDISP;
assign #(in_delay) PHYEMAC0SIGNALDET_delay = PHYEMAC0SIGNALDET;
assign #(in_delay) PHYEMAC0TXBUFERR_delay = PHYEMAC0TXBUFERR;
assign #(in_delay) PHYEMAC1COL_delay = PHYEMAC1COL;
assign #(in_delay) PHYEMAC1CRS_delay = PHYEMAC1CRS;
assign #(in_delay) PHYEMAC1MCLKIN_delay = PHYEMAC1MCLKIN;
assign #(in_delay) PHYEMAC1MDIN_delay = PHYEMAC1MDIN;
assign #(in_delay) PHYEMAC1PHYAD_delay[4:0] = PHYEMAC1PHYAD[4:0];
assign #(in_delay) PHYEMAC1RXBUFERR_delay = PHYEMAC1RXBUFERR;
assign #(in_delay) PHYEMAC1RXBUFSTATUS_delay[1:0] = PHYEMAC1RXBUFSTATUS[1:0];
assign #(in_delay) PHYEMAC1RXCHARISCOMMA_delay = PHYEMAC1RXCHARISCOMMA;
assign #(in_delay) PHYEMAC1RXCHARISK_delay = PHYEMAC1RXCHARISK;
assign #(in_delay) PHYEMAC1RXCHECKINGCRC_delay = PHYEMAC1RXCHECKINGCRC;
assign #(in_delay) PHYEMAC1RXCLKCORCNT_delay[2:0] = PHYEMAC1RXCLKCORCNT[2:0];
assign #(in_delay) PHYEMAC1RXCOMMADET_delay = PHYEMAC1RXCOMMADET;
assign #(in_delay) PHYEMAC1RXDISPERR_delay = PHYEMAC1RXDISPERR;
assign #(in_delay) PHYEMAC1RXDV_delay = PHYEMAC1RXDV;
assign #(in_delay) PHYEMAC1RXD_delay[7:0] = PHYEMAC1RXD[7:0];
assign #(in_delay) PHYEMAC1RXER_delay = PHYEMAC1RXER;
assign #(in_delay) PHYEMAC1RXLOSSOFSYNC_delay[1:0] = PHYEMAC1RXLOSSOFSYNC[1:0];
assign #(in_delay) PHYEMAC1RXNOTINTABLE_delay = PHYEMAC1RXNOTINTABLE;
assign #(in_delay) PHYEMAC1RXRUNDISP_delay = PHYEMAC1RXRUNDISP;
assign #(in_delay) PHYEMAC1SIGNALDET_delay = PHYEMAC1SIGNALDET;
assign #(in_delay) PHYEMAC1TXBUFERR_delay = PHYEMAC1TXBUFERR;
assign #(in_delay) RESET_delay = RESET;
assign #(in_delay) TIEEMAC0CONFIGVEC_delay[79:0] = TIEEMAC0CONFIGVEC[79:0];
assign #(in_delay) TIEEMAC0UNICASTADDR_delay[47:0] = TIEEMAC0UNICASTADDR[47:0];
assign #(in_delay) TIEEMAC1CONFIGVEC_delay[79:0] = TIEEMAC1CONFIGVEC[79:0];
assign #(in_delay) TIEEMAC1UNICASTADDR_delay[47:0] = TIEEMAC1UNICASTADDR[47:0];
assign #(out_delay) DCRHOSTDONEIR = DCRHOSTDONEIR_delay;
assign #(out_delay) EMAC0CLIENTANINTERRUPT = EMAC0CLIENTANINTERRUPT_delay;
assign #(out_delay) EMAC0CLIENTRXBADFRAME = EMAC0CLIENTRXBADFRAME_delay;
assign #(out_delay) EMAC0CLIENTRXDVLD = EMAC0CLIENTRXDVLD_delay;
assign #(out_delay) EMAC0CLIENTRXDVLDMSW = EMAC0CLIENTRXDVLDMSW_delay;
assign #(out_delay) EMAC0CLIENTRXDVREG6 = EMAC0CLIENTRXDVREG6_delay;
assign #(out_delay) EMAC0CLIENTRXD[15:0] = EMAC0CLIENTRXD_delay[15:0];
assign #(out_delay) EMAC0CLIENTRXFRAMEDROP = EMAC0CLIENTRXFRAMEDROP_delay;
assign #(out_delay) EMAC0CLIENTRXGOODFRAME = EMAC0CLIENTRXGOODFRAME_delay;
assign #(out_delay) EMAC0CLIENTRXSTATSBYTEVLD = EMAC0CLIENTRXSTATSBYTEVLD_delay;
assign #(out_delay) EMAC0CLIENTRXSTATSVLD = EMAC0CLIENTRXSTATSVLD_delay;
assign #(out_delay) EMAC0CLIENTRXSTATS[6:0] = EMAC0CLIENTRXSTATS_delay[6:0];
assign #(out_delay) EMAC0CLIENTTXACK = EMAC0CLIENTTXACK_delay;
assign #(out_delay) EMAC0CLIENTTXCOLLISION = EMAC0CLIENTTXCOLLISION_delay;
assign #(out_delay) EMAC0CLIENTTXRETRANSMIT = EMAC0CLIENTTXRETRANSMIT_delay;
assign #(out_delay) EMAC0CLIENTTXSTATS = EMAC0CLIENTTXSTATS_delay;
assign #(out_delay) EMAC0CLIENTTXSTATSBYTEVLD = EMAC0CLIENTTXSTATSBYTEVLD_delay;
assign #(out_delay) EMAC0CLIENTTXSTATSVLD = EMAC0CLIENTTXSTATSVLD_delay;
assign #(out_delay) EMAC0PHYENCOMMAALIGN = EMAC0PHYENCOMMAALIGN_delay;
assign #(out_delay) EMAC0PHYLOOPBACKMSB = EMAC0PHYLOOPBACKMSB_delay;
assign #(out_delay) EMAC0PHYMCLKOUT = EMAC0PHYMCLKOUT_delay;
assign #(out_delay) EMAC0PHYMDOUT = EMAC0PHYMDOUT_delay;
assign #(out_delay) EMAC0PHYMDTRI = EMAC0PHYMDTRI_delay;
assign #(out_delay) EMAC0PHYMGTRXRESET = EMAC0PHYMGTRXRESET_delay;
assign #(out_delay) EMAC0PHYMGTTXRESET = EMAC0PHYMGTTXRESET_delay;
assign #(out_delay) EMAC0PHYPOWERDOWN = EMAC0PHYPOWERDOWN_delay;
assign #(out_delay) EMAC0PHYSYNCACQSTATUS = EMAC0PHYSYNCACQSTATUS_delay;
assign #(out_delay) EMAC0PHYTXCHARDISPMODE = EMAC0PHYTXCHARDISPMODE_delay;
assign #(out_delay) EMAC0PHYTXCHARDISPVAL = EMAC0PHYTXCHARDISPVAL_delay;
assign #(out_delay) EMAC0PHYTXCHARISK = EMAC0PHYTXCHARISK_delay;
assign #(out_delay) EMAC0PHYTXD[7:0] = EMAC0PHYTXD_delay[7:0];
assign #(out_delay) EMAC0PHYTXEN = EMAC0PHYTXEN_delay;
assign #(out_delay) EMAC0PHYTXER = EMAC0PHYTXER_delay;
assign #(out_delay) EMAC1CLIENTANINTERRUPT = EMAC1CLIENTANINTERRUPT_delay;
assign #(out_delay) EMAC1CLIENTRXBADFRAME = EMAC1CLIENTRXBADFRAME_delay;
assign #(out_delay) EMAC1CLIENTRXDVLD = EMAC1CLIENTRXDVLD_delay;
assign #(out_delay) EMAC1CLIENTRXDVLDMSW = EMAC1CLIENTRXDVLDMSW_delay;
assign #(out_delay) EMAC1CLIENTRXDVREG6 = EMAC1CLIENTRXDVREG6_delay;
assign #(out_delay) EMAC1CLIENTRXD[15:0] = EMAC1CLIENTRXD_delay[15:0];
assign #(out_delay) EMAC1CLIENTRXFRAMEDROP = EMAC1CLIENTRXFRAMEDROP_delay;
assign #(out_delay) EMAC1CLIENTRXGOODFRAME = EMAC1CLIENTRXGOODFRAME_delay;
assign #(out_delay) EMAC1CLIENTRXSTATSBYTEVLD = EMAC1CLIENTRXSTATSBYTEVLD_delay;
assign #(out_delay) EMAC1CLIENTRXSTATSVLD = EMAC1CLIENTRXSTATSVLD_delay;
assign #(out_delay) EMAC1CLIENTRXSTATS[6:0] = EMAC1CLIENTRXSTATS_delay[6:0];
assign #(out_delay) EMAC1CLIENTTXACK = EMAC1CLIENTTXACK_delay;
assign #(out_delay) EMAC1CLIENTTXCOLLISION = EMAC1CLIENTTXCOLLISION_delay;
assign #(out_delay) EMAC1CLIENTTXRETRANSMIT = EMAC1CLIENTTXRETRANSMIT_delay;
assign #(out_delay) EMAC1CLIENTTXSTATS = EMAC1CLIENTTXSTATS_delay;
assign #(out_delay) EMAC1CLIENTTXSTATSBYTEVLD = EMAC1CLIENTTXSTATSBYTEVLD_delay;
assign #(out_delay) EMAC1CLIENTTXSTATSVLD = EMAC1CLIENTTXSTATSVLD_delay;
assign #(out_delay) EMAC1PHYENCOMMAALIGN = EMAC1PHYENCOMMAALIGN_delay;
assign #(out_delay) EMAC1PHYLOOPBACKMSB = EMAC1PHYLOOPBACKMSB_delay;
assign #(out_delay) EMAC1PHYMCLKOUT = EMAC1PHYMCLKOUT_delay;
assign #(out_delay) EMAC1PHYMDOUT = EMAC1PHYMDOUT_delay;
assign #(out_delay) EMAC1PHYMDTRI = EMAC1PHYMDTRI_delay;
assign #(out_delay) EMAC1PHYMGTRXRESET = EMAC1PHYMGTRXRESET_delay;
assign #(out_delay) EMAC1PHYMGTTXRESET = EMAC1PHYMGTTXRESET_delay;
assign #(out_delay) EMAC1PHYPOWERDOWN = EMAC1PHYPOWERDOWN_delay;
assign #(out_delay) EMAC1PHYSYNCACQSTATUS = EMAC1PHYSYNCACQSTATUS_delay;
assign #(out_delay) EMAC1PHYTXCHARDISPMODE = EMAC1PHYTXCHARDISPMODE_delay;
assign #(out_delay) EMAC1PHYTXCHARDISPVAL = EMAC1PHYTXCHARDISPVAL_delay;
assign #(out_delay) EMAC1PHYTXCHARISK = EMAC1PHYTXCHARISK_delay;
assign #(out_delay) EMAC1PHYTXD[7:0] = EMAC1PHYTXD_delay[7:0];
assign #(out_delay) EMAC1PHYTXEN = EMAC1PHYTXEN_delay;
assign #(out_delay) EMAC1PHYTXER = EMAC1PHYTXER_delay;
assign #(out_delay) EMACDCRACK = EMACDCRACK_delay;
assign #(out_delay) EMACDCRDBUS[0:31] = EMACDCRDBUS_delay[0:31];
assign #(out_delay) HOSTMIIMRDY = HOSTMIIMRDY_delay;
assign #(out_delay) HOSTRDDATA[31:0] = HOSTRDDATA_delay[31:0];

EMAC_SWIFT EMAC_SWIFT (
	.CLIENTEMAC0DCMLOCKED (CLIENTEMAC0DCMLOCKED_delay),
	.CLIENTEMAC0PAUSEREQ (CLIENTEMAC0PAUSEREQ_delay),
	.CLIENTEMAC0PAUSEVAL (CLIENTEMAC0PAUSEVAL_delay),
	.CLIENTEMAC0RXCLIENTCLKIN (CLIENTEMAC0RXCLIENTCLKIN),
	.CLIENTEMAC0TXCLIENTCLKIN (CLIENTEMAC0TXCLIENTCLKIN),
	.CLIENTEMAC0TXD (CLIENTEMAC0TXD_delay),
	.CLIENTEMAC0TXDVLD (CLIENTEMAC0TXDVLD_delay),
	.CLIENTEMAC0TXDVLDMSW (CLIENTEMAC0TXDVLDMSW_delay),
	.CLIENTEMAC0TXFIRSTBYTE (CLIENTEMAC0TXFIRSTBYTE_delay),
	.CLIENTEMAC0TXGMIIMIICLKIN (CLIENTEMAC0TXGMIIMIICLKIN),
	.CLIENTEMAC0TXIFGDELAY (CLIENTEMAC0TXIFGDELAY_delay),
	.CLIENTEMAC0TXUNDERRUN (CLIENTEMAC0TXUNDERRUN_delay),
	.CLIENTEMAC1DCMLOCKED (CLIENTEMAC1DCMLOCKED_delay),
	.CLIENTEMAC1PAUSEREQ (CLIENTEMAC1PAUSEREQ_delay),
	.CLIENTEMAC1PAUSEVAL (CLIENTEMAC1PAUSEVAL_delay),
	.CLIENTEMAC1RXCLIENTCLKIN (CLIENTEMAC1RXCLIENTCLKIN),
	.CLIENTEMAC1TXCLIENTCLKIN (CLIENTEMAC1TXCLIENTCLKIN),
	.CLIENTEMAC1TXD (CLIENTEMAC1TXD_delay),
	.CLIENTEMAC1TXDVLD (CLIENTEMAC1TXDVLD_delay),
	.CLIENTEMAC1TXDVLDMSW (CLIENTEMAC1TXDVLDMSW_delay),
	.CLIENTEMAC1TXFIRSTBYTE (CLIENTEMAC1TXFIRSTBYTE_delay),
	.CLIENTEMAC1TXGMIIMIICLKIN (CLIENTEMAC1TXGMIIMIICLKIN),
	.CLIENTEMAC1TXIFGDELAY (CLIENTEMAC1TXIFGDELAY_delay),
	.CLIENTEMAC1TXUNDERRUN (CLIENTEMAC1TXUNDERRUN_delay),
	.DCREMACABUS (DCREMACABUS_delay[8:9]),
	.DCREMACCLK (DCREMACCLK),
	.DCREMACDBUS (DCREMACDBUS_delay[0:31]),
	.DCREMACENABLE (DCREMACENABLE_delay),
	.DCREMACREAD (DCREMACREAD_delay),
	.DCREMACWRITE (DCREMACWRITE_delay),
	.DCRHOSTDONEIR (DCRHOSTDONEIR_delay),
	.EMAC0CLIENTANINTERRUPT (EMAC0CLIENTANINTERRUPT_delay),
	.EMAC0CLIENTRXBADFRAME (EMAC0CLIENTRXBADFRAME_delay),
	.EMAC0CLIENTRXCLIENTCLKOUT (EMAC0CLIENTRXCLIENTCLKOUT),
	.EMAC0CLIENTRXD (EMAC0CLIENTRXD_delay),
	.EMAC0CLIENTRXDVLD (EMAC0CLIENTRXDVLD_delay),
	.EMAC0CLIENTRXDVLDMSW (EMAC0CLIENTRXDVLDMSW_delay),
	.EMAC0CLIENTRXDVREG6 (EMAC0CLIENTRXDVREG6_delay),
	.EMAC0CLIENTRXFRAMEDROP (EMAC0CLIENTRXFRAMEDROP_delay),
	.EMAC0CLIENTRXGOODFRAME (EMAC0CLIENTRXGOODFRAME_delay),
	.EMAC0CLIENTRXSTATS (EMAC0CLIENTRXSTATS_delay),
	.EMAC0CLIENTRXSTATSBYTEVLD (EMAC0CLIENTRXSTATSBYTEVLD_delay),
	.EMAC0CLIENTRXSTATSVLD (EMAC0CLIENTRXSTATSVLD_delay),
	.EMAC0CLIENTTXACK (EMAC0CLIENTTXACK_delay),
	.EMAC0CLIENTTXCLIENTCLKOUT (EMAC0CLIENTTXCLIENTCLKOUT),
	.EMAC0CLIENTTXCOLLISION (EMAC0CLIENTTXCOLLISION_delay),
	.EMAC0CLIENTTXGMIIMIICLKOUT (EMAC0CLIENTTXGMIIMIICLKOUT),
	.EMAC0CLIENTTXRETRANSMIT (EMAC0CLIENTTXRETRANSMIT_delay),
	.EMAC0CLIENTTXSTATS (EMAC0CLIENTTXSTATS_delay),
	.EMAC0CLIENTTXSTATSBYTEVLD (EMAC0CLIENTTXSTATSBYTEVLD_delay),
	.EMAC0CLIENTTXSTATSVLD (EMAC0CLIENTTXSTATSVLD_delay),
	.EMAC0PHYENCOMMAALIGN (EMAC0PHYENCOMMAALIGN_delay),
	.EMAC0PHYLOOPBACKMSB (EMAC0PHYLOOPBACKMSB_delay),
	.EMAC0PHYMCLKOUT (EMAC0PHYMCLKOUT_delay),
	.EMAC0PHYMDOUT (EMAC0PHYMDOUT_delay),
	.EMAC0PHYMDTRI (EMAC0PHYMDTRI_delay),
	.EMAC0PHYMGTRXRESET (EMAC0PHYMGTRXRESET_delay),
	.EMAC0PHYMGTTXRESET (EMAC0PHYMGTTXRESET_delay),
	.EMAC0PHYPOWERDOWN (EMAC0PHYPOWERDOWN_delay),
	.EMAC0PHYSYNCACQSTATUS (EMAC0PHYSYNCACQSTATUS_delay),
	.EMAC0PHYTXCHARDISPMODE (EMAC0PHYTXCHARDISPMODE_delay),
	.EMAC0PHYTXCHARDISPVAL (EMAC0PHYTXCHARDISPVAL_delay),
	.EMAC0PHYTXCHARISK (EMAC0PHYTXCHARISK_delay),
	.EMAC0PHYTXCLK (EMAC0PHYTXCLK),
	.EMAC0PHYTXD (EMAC0PHYTXD_delay),
	.EMAC0PHYTXEN (EMAC0PHYTXEN_delay),
	.EMAC0PHYTXER (EMAC0PHYTXER_delay),
	.EMAC1CLIENTANINTERRUPT (EMAC1CLIENTANINTERRUPT_delay),
	.EMAC1CLIENTRXBADFRAME (EMAC1CLIENTRXBADFRAME_delay),
	.EMAC1CLIENTRXCLIENTCLKOUT (EMAC1CLIENTRXCLIENTCLKOUT),
	.EMAC1CLIENTRXD (EMAC1CLIENTRXD_delay),
	.EMAC1CLIENTRXDVLD (EMAC1CLIENTRXDVLD_delay),
	.EMAC1CLIENTRXDVLDMSW (EMAC1CLIENTRXDVLDMSW_delay),
	.EMAC1CLIENTRXDVREG6 (EMAC1CLIENTRXDVREG6_delay),
	.EMAC1CLIENTRXFRAMEDROP (EMAC1CLIENTRXFRAMEDROP_delay),
	.EMAC1CLIENTRXGOODFRAME (EMAC1CLIENTRXGOODFRAME_delay),
	.EMAC1CLIENTRXSTATS (EMAC1CLIENTRXSTATS_delay),
	.EMAC1CLIENTRXSTATSBYTEVLD (EMAC1CLIENTRXSTATSBYTEVLD_delay),
	.EMAC1CLIENTRXSTATSVLD (EMAC1CLIENTRXSTATSVLD_delay),
	.EMAC1CLIENTTXACK (EMAC1CLIENTTXACK_delay),
	.EMAC1CLIENTTXCLIENTCLKOUT (EMAC1CLIENTTXCLIENTCLKOUT),
	.EMAC1CLIENTTXCOLLISION (EMAC1CLIENTTXCOLLISION_delay),
	.EMAC1CLIENTTXGMIIMIICLKOUT (EMAC1CLIENTTXGMIIMIICLKOUT),
	.EMAC1CLIENTTXRETRANSMIT (EMAC1CLIENTTXRETRANSMIT_delay),
	.EMAC1CLIENTTXSTATS (EMAC1CLIENTTXSTATS_delay),
	.EMAC1CLIENTTXSTATSBYTEVLD (EMAC1CLIENTTXSTATSBYTEVLD_delay),
	.EMAC1CLIENTTXSTATSVLD (EMAC1CLIENTTXSTATSVLD_delay),
	.EMAC1PHYENCOMMAALIGN (EMAC1PHYENCOMMAALIGN_delay),
	.EMAC1PHYLOOPBACKMSB (EMAC1PHYLOOPBACKMSB_delay),
	.EMAC1PHYMCLKOUT (EMAC1PHYMCLKOUT_delay),
	.EMAC1PHYMDOUT (EMAC1PHYMDOUT_delay),
	.EMAC1PHYMDTRI (EMAC1PHYMDTRI_delay),
	.EMAC1PHYMGTRXRESET (EMAC1PHYMGTRXRESET_delay),
	.EMAC1PHYMGTTXRESET (EMAC1PHYMGTTXRESET_delay),
	.EMAC1PHYPOWERDOWN (EMAC1PHYPOWERDOWN_delay),
	.EMAC1PHYSYNCACQSTATUS (EMAC1PHYSYNCACQSTATUS_delay),
	.EMAC1PHYTXCHARDISPMODE (EMAC1PHYTXCHARDISPMODE_delay),
	.EMAC1PHYTXCHARDISPVAL (EMAC1PHYTXCHARDISPVAL_delay),
	.EMAC1PHYTXCHARISK (EMAC1PHYTXCHARISK_delay),
	.EMAC1PHYTXCLK (EMAC1PHYTXCLK),
	.EMAC1PHYTXD (EMAC1PHYTXD_delay),
	.EMAC1PHYTXEN (EMAC1PHYTXEN_delay),
	.EMAC1PHYTXER (EMAC1PHYTXER_delay),
	.EMACDCRACK (EMACDCRACK_delay),
	.EMACDCRDBUS (EMACDCRDBUS_delay[0:31]),
	.HOSTADDR (HOSTADDR_delay),
	.HOSTCLK (HOSTCLK),
	.HOSTEMAC1SEL (HOSTEMAC1SEL_delay),
	.HOSTMIIMRDY (HOSTMIIMRDY_delay),
	.HOSTMIIMSEL (HOSTMIIMSEL_delay),
	.HOSTOPCODE (HOSTOPCODE_delay),
	.HOSTRDDATA (HOSTRDDATA_delay),
	.HOSTREQ (HOSTREQ_delay),
	.HOSTWRDATA (HOSTWRDATA_delay),
	.PHYEMAC0COL (PHYEMAC0COL_delay),
	.PHYEMAC0CRS (PHYEMAC0CRS_delay),
	.PHYEMAC0GTXCLK (PHYEMAC0GTXCLK),
	.PHYEMAC0MCLKIN (PHYEMAC0MCLKIN_delay),
	.PHYEMAC0MDIN (PHYEMAC0MDIN_delay),
	.PHYEMAC0MIITXCLK (PHYEMAC0MIITXCLK),
	.PHYEMAC0PHYAD (PHYEMAC0PHYAD_delay),
	.PHYEMAC0RXBUFERR (PHYEMAC0RXBUFERR_delay),
	.PHYEMAC0RXBUFSTATUS (PHYEMAC0RXBUFSTATUS_delay),
	.PHYEMAC0RXCHARISCOMMA (PHYEMAC0RXCHARISCOMMA_delay),
	.PHYEMAC0RXCHARISK (PHYEMAC0RXCHARISK_delay),
	.PHYEMAC0RXCHECKINGCRC (PHYEMAC0RXCHECKINGCRC_delay),
	.PHYEMAC0RXCLK (PHYEMAC0RXCLK),
	.PHYEMAC0RXCLKCORCNT (PHYEMAC0RXCLKCORCNT_delay),
	.PHYEMAC0RXCOMMADET (PHYEMAC0RXCOMMADET_delay),
	.PHYEMAC0RXD (PHYEMAC0RXD_delay),
	.PHYEMAC0RXDISPERR (PHYEMAC0RXDISPERR_delay),
	.PHYEMAC0RXDV (PHYEMAC0RXDV_delay),
	.PHYEMAC0RXER (PHYEMAC0RXER_delay),
	.PHYEMAC0RXLOSSOFSYNC (PHYEMAC0RXLOSSOFSYNC_delay),
	.PHYEMAC0RXNOTINTABLE (PHYEMAC0RXNOTINTABLE_delay),
	.PHYEMAC0RXRUNDISP (PHYEMAC0RXRUNDISP_delay),
	.PHYEMAC0SIGNALDET (PHYEMAC0SIGNALDET_delay),
	.PHYEMAC0TXBUFERR (PHYEMAC0TXBUFERR_delay),
	.PHYEMAC1COL (PHYEMAC1COL_delay),
	.PHYEMAC1CRS (PHYEMAC1CRS_delay), 
	.PHYEMAC1GTXCLK (PHYEMAC1GTXCLK),
	.PHYEMAC1MCLKIN (PHYEMAC1MCLKIN_delay),
	.PHYEMAC1MDIN (PHYEMAC1MDIN_delay),
	.PHYEMAC1MIITXCLK (PHYEMAC1MIITXCLK),
	.PHYEMAC1PHYAD (PHYEMAC1PHYAD_delay),
	.PHYEMAC1RXBUFERR (PHYEMAC1RXBUFERR_delay),
	.PHYEMAC1RXBUFSTATUS (PHYEMAC1RXBUFSTATUS_delay),
	.PHYEMAC1RXCHARISCOMMA (PHYEMAC1RXCHARISCOMMA_delay),
	.PHYEMAC1RXCHARISK (PHYEMAC1RXCHARISK_delay),
	.PHYEMAC1RXCHECKINGCRC (PHYEMAC1RXCHECKINGCRC_delay),
	.PHYEMAC1RXCLK (PHYEMAC1RXCLK),
	.PHYEMAC1RXCLKCORCNT (PHYEMAC1RXCLKCORCNT_delay),
	.PHYEMAC1RXCOMMADET (PHYEMAC1RXCOMMADET_delay),
	.PHYEMAC1RXD (PHYEMAC1RXD_delay),
	.PHYEMAC1RXDISPERR (PHYEMAC1RXDISPERR_delay),
	.PHYEMAC1RXDV (PHYEMAC1RXDV_delay),
	.PHYEMAC1RXER (PHYEMAC1RXER_delay),
	.PHYEMAC1RXLOSSOFSYNC (PHYEMAC1RXLOSSOFSYNC_delay),
	.PHYEMAC1RXNOTINTABLE (PHYEMAC1RXNOTINTABLE_delay),
	.PHYEMAC1RXRUNDISP (PHYEMAC1RXRUNDISP_delay),
	.PHYEMAC1SIGNALDET (PHYEMAC1SIGNALDET_delay),
	.PHYEMAC1TXBUFERR (PHYEMAC1TXBUFERR_delay),
	.RESET (RESET_delay),
	.TIEEMAC0CONFIGVEC (TIEEMAC0CONFIGVEC_delay),
	.TIEEMAC0UNICASTADDR (TIEEMAC0UNICASTADDR_delay),
	.TIEEMAC1CONFIGVEC (TIEEMAC1CONFIGVEC_delay),
	.TIEEMAC1UNICASTADDR (TIEEMAC1UNICASTADDR_delay)
);

endmodule
