// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/GND.v,v 1.8.22.1 2003/11/18 20:41:34 wloo Exp $

/*

FUNCTION	: GND cell

*/

`timescale  100 ps / 10 ps


module GND(G);

    output G;

	assign G = 1'b0;

endmodule

