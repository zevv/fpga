// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/CAPTURE_SPARTAN2.v,v 1.8.22.1 2003/11/18 20:41:33 wloo Exp $
/*

FUNCTION	: Special Function Cell, CAPTURE_SPARTAN2

*/

`timescale  100 ps / 10 ps


module CAPTURE_SPARTAN2 (CAP, CLK);

    input  CAP, CLK;

endmodule

