// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/CAPTURE_VIRTEX4.v,v 1.1.6.6 2004/05/12 19:07:22 patrickp Exp $
/*

FUNCTION	: Special Function Cell, CAPTURE_VIRTEX4

*/

`timescale  100 ps / 10 ps


module CAPTURE_VIRTEX4 (CAP, CLK);

    input  CAP, CLK;

    parameter ONESHOT = "TRUE";
    
endmodule
